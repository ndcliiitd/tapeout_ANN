VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1209.080 200.000 1209.680 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1375.000 200.000 1375.600 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1540.920 200.000 1541.520 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1706.840 200.000 1707.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1872.760 200.000 1873.360 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2038.680 200.000 2039.280 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2204.600 200.000 2205.200 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2370.520 200.000 2371.120 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2536.440 200.000 2537.040 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2702.360 200.000 2702.960 ;
    END
  END io_in[19]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2868.280 200.000 2868.880 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2934.920 4.000 2935.520 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2760.840 4.000 2761.440 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2586.760 4.000 2587.360 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2412.680 4.000 2413.280 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2238.600 4.000 2239.200 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2064.520 4.000 2065.120 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1890.440 4.000 1891.040 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1716.360 4.000 1716.960 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1542.280 4.000 1542.880 ;
    END
  END io_in[29]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1368.200 4.000 1368.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_in[37]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 711.320 200.000 711.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 877.240 200.000 877.840 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1043.160 200.000 1043.760 ;
    END
  END io_in[9]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1292.040 200.000 1292.640 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1457.960 200.000 1458.560 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1623.880 200.000 1624.480 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1789.800 200.000 1790.400 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1955.720 200.000 1956.320 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2121.640 200.000 2122.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2287.560 200.000 2288.160 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2453.480 200.000 2454.080 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2619.400 200.000 2620.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2785.320 200.000 2785.920 ;
    END
  END io_oeb[19]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2951.240 200.000 2951.840 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2847.880 4.000 2848.480 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2673.800 4.000 2674.400 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2499.720 4.000 2500.320 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2325.640 4.000 2326.240 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2151.560 4.000 2152.160 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1977.480 4.000 1978.080 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1803.400 4.000 1804.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1629.320 4.000 1629.920 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.160 4.000 1281.760 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1107.080 4.000 1107.680 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 130.600 200.000 131.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 296.520 200.000 297.120 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 462.440 200.000 463.040 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 628.360 200.000 628.960 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 794.280 200.000 794.880 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 960.200 200.000 960.800 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1126.120 200.000 1126.720 ;
    END
  END io_oeb[9]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 47.640 200.000 48.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 213.560 200.000 214.160 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 379.480 200.000 380.080 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 545.400 200.000 546.000 ;
    END
  END io_out[6]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 195.430 2986.800 ;
      LAYER met2 ;
        RECT 4.690 4.280 195.400 2986.745 ;
        RECT 4.690 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 195.400 4.280 ;
      LAYER met3 ;
        RECT 3.990 2952.240 196.000 2986.725 ;
        RECT 3.990 2950.840 195.600 2952.240 ;
        RECT 3.990 2935.920 196.000 2950.840 ;
        RECT 4.400 2934.520 196.000 2935.920 ;
        RECT 3.990 2869.280 196.000 2934.520 ;
        RECT 3.990 2867.880 195.600 2869.280 ;
        RECT 3.990 2848.880 196.000 2867.880 ;
        RECT 4.400 2847.480 196.000 2848.880 ;
        RECT 3.990 2786.320 196.000 2847.480 ;
        RECT 3.990 2784.920 195.600 2786.320 ;
        RECT 3.990 2761.840 196.000 2784.920 ;
        RECT 4.400 2760.440 196.000 2761.840 ;
        RECT 3.990 2703.360 196.000 2760.440 ;
        RECT 3.990 2701.960 195.600 2703.360 ;
        RECT 3.990 2674.800 196.000 2701.960 ;
        RECT 4.400 2673.400 196.000 2674.800 ;
        RECT 3.990 2620.400 196.000 2673.400 ;
        RECT 3.990 2619.000 195.600 2620.400 ;
        RECT 3.990 2587.760 196.000 2619.000 ;
        RECT 4.400 2586.360 196.000 2587.760 ;
        RECT 3.990 2537.440 196.000 2586.360 ;
        RECT 3.990 2536.040 195.600 2537.440 ;
        RECT 3.990 2500.720 196.000 2536.040 ;
        RECT 4.400 2499.320 196.000 2500.720 ;
        RECT 3.990 2454.480 196.000 2499.320 ;
        RECT 3.990 2453.080 195.600 2454.480 ;
        RECT 3.990 2413.680 196.000 2453.080 ;
        RECT 4.400 2412.280 196.000 2413.680 ;
        RECT 3.990 2371.520 196.000 2412.280 ;
        RECT 3.990 2370.120 195.600 2371.520 ;
        RECT 3.990 2326.640 196.000 2370.120 ;
        RECT 4.400 2325.240 196.000 2326.640 ;
        RECT 3.990 2288.560 196.000 2325.240 ;
        RECT 3.990 2287.160 195.600 2288.560 ;
        RECT 3.990 2239.600 196.000 2287.160 ;
        RECT 4.400 2238.200 196.000 2239.600 ;
        RECT 3.990 2205.600 196.000 2238.200 ;
        RECT 3.990 2204.200 195.600 2205.600 ;
        RECT 3.990 2152.560 196.000 2204.200 ;
        RECT 4.400 2151.160 196.000 2152.560 ;
        RECT 3.990 2122.640 196.000 2151.160 ;
        RECT 3.990 2121.240 195.600 2122.640 ;
        RECT 3.990 2065.520 196.000 2121.240 ;
        RECT 4.400 2064.120 196.000 2065.520 ;
        RECT 3.990 2039.680 196.000 2064.120 ;
        RECT 3.990 2038.280 195.600 2039.680 ;
        RECT 3.990 1978.480 196.000 2038.280 ;
        RECT 4.400 1977.080 196.000 1978.480 ;
        RECT 3.990 1956.720 196.000 1977.080 ;
        RECT 3.990 1955.320 195.600 1956.720 ;
        RECT 3.990 1891.440 196.000 1955.320 ;
        RECT 4.400 1890.040 196.000 1891.440 ;
        RECT 3.990 1873.760 196.000 1890.040 ;
        RECT 3.990 1872.360 195.600 1873.760 ;
        RECT 3.990 1804.400 196.000 1872.360 ;
        RECT 4.400 1803.000 196.000 1804.400 ;
        RECT 3.990 1790.800 196.000 1803.000 ;
        RECT 3.990 1789.400 195.600 1790.800 ;
        RECT 3.990 1717.360 196.000 1789.400 ;
        RECT 4.400 1715.960 196.000 1717.360 ;
        RECT 3.990 1707.840 196.000 1715.960 ;
        RECT 3.990 1706.440 195.600 1707.840 ;
        RECT 3.990 1630.320 196.000 1706.440 ;
        RECT 4.400 1628.920 196.000 1630.320 ;
        RECT 3.990 1624.880 196.000 1628.920 ;
        RECT 3.990 1623.480 195.600 1624.880 ;
        RECT 3.990 1543.280 196.000 1623.480 ;
        RECT 4.400 1541.920 196.000 1543.280 ;
        RECT 4.400 1541.880 195.600 1541.920 ;
        RECT 3.990 1540.520 195.600 1541.880 ;
        RECT 3.990 1458.960 196.000 1540.520 ;
        RECT 3.990 1457.560 195.600 1458.960 ;
        RECT 3.990 1456.240 196.000 1457.560 ;
        RECT 4.400 1454.840 196.000 1456.240 ;
        RECT 3.990 1376.000 196.000 1454.840 ;
        RECT 3.990 1374.600 195.600 1376.000 ;
        RECT 3.990 1369.200 196.000 1374.600 ;
        RECT 4.400 1367.800 196.000 1369.200 ;
        RECT 3.990 1293.040 196.000 1367.800 ;
        RECT 3.990 1291.640 195.600 1293.040 ;
        RECT 3.990 1282.160 196.000 1291.640 ;
        RECT 4.400 1280.760 196.000 1282.160 ;
        RECT 3.990 1210.080 196.000 1280.760 ;
        RECT 3.990 1208.680 195.600 1210.080 ;
        RECT 3.990 1195.120 196.000 1208.680 ;
        RECT 4.400 1193.720 196.000 1195.120 ;
        RECT 3.990 1127.120 196.000 1193.720 ;
        RECT 3.990 1125.720 195.600 1127.120 ;
        RECT 3.990 1108.080 196.000 1125.720 ;
        RECT 4.400 1106.680 196.000 1108.080 ;
        RECT 3.990 1044.160 196.000 1106.680 ;
        RECT 3.990 1042.760 195.600 1044.160 ;
        RECT 3.990 1021.040 196.000 1042.760 ;
        RECT 4.400 1019.640 196.000 1021.040 ;
        RECT 3.990 961.200 196.000 1019.640 ;
        RECT 3.990 959.800 195.600 961.200 ;
        RECT 3.990 934.000 196.000 959.800 ;
        RECT 4.400 932.600 196.000 934.000 ;
        RECT 3.990 878.240 196.000 932.600 ;
        RECT 3.990 876.840 195.600 878.240 ;
        RECT 3.990 846.960 196.000 876.840 ;
        RECT 4.400 845.560 196.000 846.960 ;
        RECT 3.990 795.280 196.000 845.560 ;
        RECT 3.990 793.880 195.600 795.280 ;
        RECT 3.990 759.920 196.000 793.880 ;
        RECT 4.400 758.520 196.000 759.920 ;
        RECT 3.990 712.320 196.000 758.520 ;
        RECT 3.990 710.920 195.600 712.320 ;
        RECT 3.990 672.880 196.000 710.920 ;
        RECT 4.400 671.480 196.000 672.880 ;
        RECT 3.990 629.360 196.000 671.480 ;
        RECT 3.990 627.960 195.600 629.360 ;
        RECT 3.990 585.840 196.000 627.960 ;
        RECT 4.400 584.440 196.000 585.840 ;
        RECT 3.990 546.400 196.000 584.440 ;
        RECT 3.990 545.000 195.600 546.400 ;
        RECT 3.990 498.800 196.000 545.000 ;
        RECT 4.400 497.400 196.000 498.800 ;
        RECT 3.990 463.440 196.000 497.400 ;
        RECT 3.990 462.040 195.600 463.440 ;
        RECT 3.990 411.760 196.000 462.040 ;
        RECT 4.400 410.360 196.000 411.760 ;
        RECT 3.990 380.480 196.000 410.360 ;
        RECT 3.990 379.080 195.600 380.480 ;
        RECT 3.990 324.720 196.000 379.080 ;
        RECT 4.400 323.320 196.000 324.720 ;
        RECT 3.990 297.520 196.000 323.320 ;
        RECT 3.990 296.120 195.600 297.520 ;
        RECT 3.990 237.680 196.000 296.120 ;
        RECT 4.400 236.280 196.000 237.680 ;
        RECT 3.990 214.560 196.000 236.280 ;
        RECT 3.990 213.160 195.600 214.560 ;
        RECT 3.990 150.640 196.000 213.160 ;
        RECT 4.400 149.240 196.000 150.640 ;
        RECT 3.990 131.600 196.000 149.240 ;
        RECT 3.990 130.200 195.600 131.600 ;
        RECT 3.990 63.600 196.000 130.200 ;
        RECT 4.400 62.200 196.000 63.600 ;
        RECT 3.990 48.640 196.000 62.200 ;
        RECT 3.990 47.240 195.600 48.640 ;
        RECT 3.990 10.715 196.000 47.240 ;
      LAYER met4 ;
        RECT 8.575 385.735 20.640 2190.785 ;
        RECT 23.040 385.735 97.440 2190.785 ;
        RECT 99.840 385.735 174.240 2190.785 ;
        RECT 176.640 385.735 183.705 2190.785 ;
  END
END user_proj_example
END LIBRARY

