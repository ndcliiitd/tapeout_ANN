// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:7] io_in;
 output [37:3] io_oeb;
 output [6:3] io_out;

 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net224;
 wire net225;
 wire net226;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire \ann.ReLU_out[0][0] ;
 wire \ann.ReLU_out[0][10] ;
 wire \ann.ReLU_out[0][11] ;
 wire \ann.ReLU_out[0][12] ;
 wire \ann.ReLU_out[0][13] ;
 wire \ann.ReLU_out[0][14] ;
 wire \ann.ReLU_out[0][15] ;
 wire \ann.ReLU_out[0][16] ;
 wire \ann.ReLU_out[0][17] ;
 wire \ann.ReLU_out[0][18] ;
 wire \ann.ReLU_out[0][19] ;
 wire \ann.ReLU_out[0][1] ;
 wire \ann.ReLU_out[0][20] ;
 wire \ann.ReLU_out[0][21] ;
 wire \ann.ReLU_out[0][22] ;
 wire \ann.ReLU_out[0][23] ;
 wire \ann.ReLU_out[0][24] ;
 wire \ann.ReLU_out[0][25] ;
 wire \ann.ReLU_out[0][26] ;
 wire \ann.ReLU_out[0][27] ;
 wire \ann.ReLU_out[0][28] ;
 wire \ann.ReLU_out[0][29] ;
 wire \ann.ReLU_out[0][2] ;
 wire \ann.ReLU_out[0][30] ;
 wire \ann.ReLU_out[0][3] ;
 wire \ann.ReLU_out[0][4] ;
 wire \ann.ReLU_out[0][5] ;
 wire \ann.ReLU_out[0][6] ;
 wire \ann.ReLU_out[0][7] ;
 wire \ann.ReLU_out[0][8] ;
 wire \ann.ReLU_out[0][9] ;
 wire \ann.ReLU_out[1][0] ;
 wire \ann.ReLU_out[1][10] ;
 wire \ann.ReLU_out[1][11] ;
 wire \ann.ReLU_out[1][12] ;
 wire \ann.ReLU_out[1][13] ;
 wire \ann.ReLU_out[1][14] ;
 wire \ann.ReLU_out[1][15] ;
 wire \ann.ReLU_out[1][16] ;
 wire \ann.ReLU_out[1][17] ;
 wire \ann.ReLU_out[1][18] ;
 wire \ann.ReLU_out[1][19] ;
 wire \ann.ReLU_out[1][1] ;
 wire \ann.ReLU_out[1][20] ;
 wire \ann.ReLU_out[1][21] ;
 wire \ann.ReLU_out[1][22] ;
 wire \ann.ReLU_out[1][23] ;
 wire \ann.ReLU_out[1][24] ;
 wire \ann.ReLU_out[1][25] ;
 wire \ann.ReLU_out[1][26] ;
 wire \ann.ReLU_out[1][27] ;
 wire \ann.ReLU_out[1][28] ;
 wire \ann.ReLU_out[1][29] ;
 wire \ann.ReLU_out[1][2] ;
 wire \ann.ReLU_out[1][30] ;
 wire \ann.ReLU_out[1][3] ;
 wire \ann.ReLU_out[1][4] ;
 wire \ann.ReLU_out[1][5] ;
 wire \ann.ReLU_out[1][6] ;
 wire \ann.ReLU_out[1][7] ;
 wire \ann.ReLU_out[1][8] ;
 wire \ann.ReLU_out[1][9] ;
 wire \ann.ReLU_out[2][0] ;
 wire \ann.ReLU_out[2][10] ;
 wire \ann.ReLU_out[2][11] ;
 wire \ann.ReLU_out[2][12] ;
 wire \ann.ReLU_out[2][13] ;
 wire \ann.ReLU_out[2][14] ;
 wire \ann.ReLU_out[2][15] ;
 wire \ann.ReLU_out[2][16] ;
 wire \ann.ReLU_out[2][17] ;
 wire \ann.ReLU_out[2][18] ;
 wire \ann.ReLU_out[2][19] ;
 wire \ann.ReLU_out[2][1] ;
 wire \ann.ReLU_out[2][20] ;
 wire \ann.ReLU_out[2][21] ;
 wire \ann.ReLU_out[2][22] ;
 wire \ann.ReLU_out[2][23] ;
 wire \ann.ReLU_out[2][24] ;
 wire \ann.ReLU_out[2][25] ;
 wire \ann.ReLU_out[2][26] ;
 wire \ann.ReLU_out[2][27] ;
 wire \ann.ReLU_out[2][28] ;
 wire \ann.ReLU_out[2][29] ;
 wire \ann.ReLU_out[2][2] ;
 wire \ann.ReLU_out[2][30] ;
 wire \ann.ReLU_out[2][3] ;
 wire \ann.ReLU_out[2][4] ;
 wire \ann.ReLU_out[2][5] ;
 wire \ann.ReLU_out[2][6] ;
 wire \ann.ReLU_out[2][7] ;
 wire \ann.ReLU_out[2][8] ;
 wire \ann.ReLU_out[2][9] ;
 wire \ann.ReLU_out[3][0] ;
 wire \ann.ReLU_out[3][10] ;
 wire \ann.ReLU_out[3][11] ;
 wire \ann.ReLU_out[3][12] ;
 wire \ann.ReLU_out[3][13] ;
 wire \ann.ReLU_out[3][14] ;
 wire \ann.ReLU_out[3][15] ;
 wire \ann.ReLU_out[3][16] ;
 wire \ann.ReLU_out[3][17] ;
 wire \ann.ReLU_out[3][18] ;
 wire \ann.ReLU_out[3][19] ;
 wire \ann.ReLU_out[3][1] ;
 wire \ann.ReLU_out[3][20] ;
 wire \ann.ReLU_out[3][21] ;
 wire \ann.ReLU_out[3][22] ;
 wire \ann.ReLU_out[3][23] ;
 wire \ann.ReLU_out[3][24] ;
 wire \ann.ReLU_out[3][25] ;
 wire \ann.ReLU_out[3][26] ;
 wire \ann.ReLU_out[3][27] ;
 wire \ann.ReLU_out[3][28] ;
 wire \ann.ReLU_out[3][29] ;
 wire \ann.ReLU_out[3][2] ;
 wire \ann.ReLU_out[3][30] ;
 wire \ann.ReLU_out[3][3] ;
 wire \ann.ReLU_out[3][4] ;
 wire \ann.ReLU_out[3][5] ;
 wire \ann.ReLU_out[3][6] ;
 wire \ann.ReLU_out[3][7] ;
 wire \ann.ReLU_out[3][8] ;
 wire \ann.ReLU_out[3][9] ;
 wire \ann.ReLU_out[4][0] ;
 wire \ann.ReLU_out[4][10] ;
 wire \ann.ReLU_out[4][11] ;
 wire \ann.ReLU_out[4][12] ;
 wire \ann.ReLU_out[4][13] ;
 wire \ann.ReLU_out[4][14] ;
 wire \ann.ReLU_out[4][15] ;
 wire \ann.ReLU_out[4][16] ;
 wire \ann.ReLU_out[4][17] ;
 wire \ann.ReLU_out[4][18] ;
 wire \ann.ReLU_out[4][19] ;
 wire \ann.ReLU_out[4][1] ;
 wire \ann.ReLU_out[4][20] ;
 wire \ann.ReLU_out[4][21] ;
 wire \ann.ReLU_out[4][22] ;
 wire \ann.ReLU_out[4][23] ;
 wire \ann.ReLU_out[4][24] ;
 wire \ann.ReLU_out[4][25] ;
 wire \ann.ReLU_out[4][26] ;
 wire \ann.ReLU_out[4][27] ;
 wire \ann.ReLU_out[4][28] ;
 wire \ann.ReLU_out[4][29] ;
 wire \ann.ReLU_out[4][2] ;
 wire \ann.ReLU_out[4][30] ;
 wire \ann.ReLU_out[4][3] ;
 wire \ann.ReLU_out[4][4] ;
 wire \ann.ReLU_out[4][5] ;
 wire \ann.ReLU_out[4][6] ;
 wire \ann.ReLU_out[4][7] ;
 wire \ann.ReLU_out[4][8] ;
 wire \ann.ReLU_out[4][9] ;
 wire \ann.ReLU_out[5][0] ;
 wire \ann.ReLU_out[5][10] ;
 wire \ann.ReLU_out[5][11] ;
 wire \ann.ReLU_out[5][12] ;
 wire \ann.ReLU_out[5][13] ;
 wire \ann.ReLU_out[5][14] ;
 wire \ann.ReLU_out[5][15] ;
 wire \ann.ReLU_out[5][16] ;
 wire \ann.ReLU_out[5][17] ;
 wire \ann.ReLU_out[5][18] ;
 wire \ann.ReLU_out[5][19] ;
 wire \ann.ReLU_out[5][1] ;
 wire \ann.ReLU_out[5][20] ;
 wire \ann.ReLU_out[5][21] ;
 wire \ann.ReLU_out[5][22] ;
 wire \ann.ReLU_out[5][23] ;
 wire \ann.ReLU_out[5][24] ;
 wire \ann.ReLU_out[5][25] ;
 wire \ann.ReLU_out[5][26] ;
 wire \ann.ReLU_out[5][27] ;
 wire \ann.ReLU_out[5][28] ;
 wire \ann.ReLU_out[5][29] ;
 wire \ann.ReLU_out[5][2] ;
 wire \ann.ReLU_out[5][30] ;
 wire \ann.ReLU_out[5][3] ;
 wire \ann.ReLU_out[5][4] ;
 wire \ann.ReLU_out[5][5] ;
 wire \ann.ReLU_out[5][6] ;
 wire \ann.ReLU_out[5][7] ;
 wire \ann.ReLU_out[5][8] ;
 wire \ann.ReLU_out[5][9] ;
 wire \ann.ReLU_out[6][0] ;
 wire \ann.ReLU_out[6][10] ;
 wire \ann.ReLU_out[6][11] ;
 wire \ann.ReLU_out[6][12] ;
 wire \ann.ReLU_out[6][13] ;
 wire \ann.ReLU_out[6][14] ;
 wire \ann.ReLU_out[6][15] ;
 wire \ann.ReLU_out[6][16] ;
 wire \ann.ReLU_out[6][17] ;
 wire \ann.ReLU_out[6][18] ;
 wire \ann.ReLU_out[6][19] ;
 wire \ann.ReLU_out[6][1] ;
 wire \ann.ReLU_out[6][20] ;
 wire \ann.ReLU_out[6][21] ;
 wire \ann.ReLU_out[6][22] ;
 wire \ann.ReLU_out[6][23] ;
 wire \ann.ReLU_out[6][24] ;
 wire \ann.ReLU_out[6][25] ;
 wire \ann.ReLU_out[6][26] ;
 wire \ann.ReLU_out[6][27] ;
 wire \ann.ReLU_out[6][28] ;
 wire \ann.ReLU_out[6][29] ;
 wire \ann.ReLU_out[6][2] ;
 wire \ann.ReLU_out[6][30] ;
 wire \ann.ReLU_out[6][3] ;
 wire \ann.ReLU_out[6][4] ;
 wire \ann.ReLU_out[6][5] ;
 wire \ann.ReLU_out[6][6] ;
 wire \ann.ReLU_out[6][7] ;
 wire \ann.ReLU_out[6][8] ;
 wire \ann.ReLU_out[6][9] ;
 wire \ann.ReLU_out[7][0] ;
 wire \ann.ReLU_out[7][10] ;
 wire \ann.ReLU_out[7][11] ;
 wire \ann.ReLU_out[7][12] ;
 wire \ann.ReLU_out[7][13] ;
 wire \ann.ReLU_out[7][14] ;
 wire \ann.ReLU_out[7][15] ;
 wire \ann.ReLU_out[7][16] ;
 wire \ann.ReLU_out[7][17] ;
 wire \ann.ReLU_out[7][18] ;
 wire \ann.ReLU_out[7][19] ;
 wire \ann.ReLU_out[7][1] ;
 wire \ann.ReLU_out[7][20] ;
 wire \ann.ReLU_out[7][21] ;
 wire \ann.ReLU_out[7][22] ;
 wire \ann.ReLU_out[7][23] ;
 wire \ann.ReLU_out[7][24] ;
 wire \ann.ReLU_out[7][25] ;
 wire \ann.ReLU_out[7][26] ;
 wire \ann.ReLU_out[7][27] ;
 wire \ann.ReLU_out[7][28] ;
 wire \ann.ReLU_out[7][29] ;
 wire \ann.ReLU_out[7][2] ;
 wire \ann.ReLU_out[7][30] ;
 wire \ann.ReLU_out[7][3] ;
 wire \ann.ReLU_out[7][4] ;
 wire \ann.ReLU_out[7][5] ;
 wire \ann.ReLU_out[7][6] ;
 wire \ann.ReLU_out[7][7] ;
 wire \ann.ReLU_out[7][8] ;
 wire \ann.ReLU_out[7][9] ;
 wire \ann.ReLU_out[8][0] ;
 wire \ann.ReLU_out[8][10] ;
 wire \ann.ReLU_out[8][11] ;
 wire \ann.ReLU_out[8][12] ;
 wire \ann.ReLU_out[8][13] ;
 wire \ann.ReLU_out[8][14] ;
 wire \ann.ReLU_out[8][15] ;
 wire \ann.ReLU_out[8][16] ;
 wire \ann.ReLU_out[8][17] ;
 wire \ann.ReLU_out[8][18] ;
 wire \ann.ReLU_out[8][19] ;
 wire \ann.ReLU_out[8][1] ;
 wire \ann.ReLU_out[8][20] ;
 wire \ann.ReLU_out[8][21] ;
 wire \ann.ReLU_out[8][22] ;
 wire \ann.ReLU_out[8][23] ;
 wire \ann.ReLU_out[8][24] ;
 wire \ann.ReLU_out[8][25] ;
 wire \ann.ReLU_out[8][26] ;
 wire \ann.ReLU_out[8][27] ;
 wire \ann.ReLU_out[8][28] ;
 wire \ann.ReLU_out[8][29] ;
 wire \ann.ReLU_out[8][2] ;
 wire \ann.ReLU_out[8][30] ;
 wire \ann.ReLU_out[8][3] ;
 wire \ann.ReLU_out[8][4] ;
 wire \ann.ReLU_out[8][5] ;
 wire \ann.ReLU_out[8][6] ;
 wire \ann.ReLU_out[8][7] ;
 wire \ann.ReLU_out[8][8] ;
 wire \ann.ReLU_out[8][9] ;
 wire \ann.ReLU_out[9][0] ;
 wire \ann.ReLU_out[9][10] ;
 wire \ann.ReLU_out[9][11] ;
 wire \ann.ReLU_out[9][12] ;
 wire \ann.ReLU_out[9][13] ;
 wire \ann.ReLU_out[9][14] ;
 wire \ann.ReLU_out[9][15] ;
 wire \ann.ReLU_out[9][16] ;
 wire \ann.ReLU_out[9][17] ;
 wire \ann.ReLU_out[9][18] ;
 wire \ann.ReLU_out[9][19] ;
 wire \ann.ReLU_out[9][1] ;
 wire \ann.ReLU_out[9][20] ;
 wire \ann.ReLU_out[9][21] ;
 wire \ann.ReLU_out[9][22] ;
 wire \ann.ReLU_out[9][23] ;
 wire \ann.ReLU_out[9][24] ;
 wire \ann.ReLU_out[9][25] ;
 wire \ann.ReLU_out[9][26] ;
 wire \ann.ReLU_out[9][27] ;
 wire \ann.ReLU_out[9][28] ;
 wire \ann.ReLU_out[9][29] ;
 wire \ann.ReLU_out[9][2] ;
 wire \ann.ReLU_out[9][30] ;
 wire \ann.ReLU_out[9][3] ;
 wire \ann.ReLU_out[9][4] ;
 wire \ann.ReLU_out[9][5] ;
 wire \ann.ReLU_out[9][6] ;
 wire \ann.ReLU_out[9][7] ;
 wire \ann.ReLU_out[9][8] ;
 wire \ann.ReLU_out[9][9] ;
 wire \ann.X[0] ;
 wire \ann.X[10] ;
 wire \ann.X[11] ;
 wire \ann.X[12] ;
 wire \ann.X[13] ;
 wire \ann.X[14] ;
 wire \ann.X[15] ;
 wire \ann.X[16] ;
 wire \ann.X[17] ;
 wire \ann.X[18] ;
 wire \ann.X[19] ;
 wire \ann.X[1] ;
 wire \ann.X[20] ;
 wire \ann.X[21] ;
 wire \ann.X[22] ;
 wire \ann.X[23] ;
 wire \ann.X[24] ;
 wire \ann.X[25] ;
 wire \ann.X[26] ;
 wire \ann.X[27] ;
 wire \ann.X[28] ;
 wire \ann.X[29] ;
 wire \ann.X[2] ;
 wire \ann.X[30] ;
 wire \ann.X[31] ;
 wire \ann.X[3] ;
 wire \ann.X[4] ;
 wire \ann.X[5] ;
 wire \ann.X[6] ;
 wire \ann.X[7] ;
 wire \ann.X[8] ;
 wire \ann.X[9] ;
 wire \ann.add_enable ;
 wire \ann.bias[0] ;
 wire \ann.bias[10] ;
 wire \ann.bias[11] ;
 wire \ann.bias[12] ;
 wire \ann.bias[13] ;
 wire \ann.bias[14] ;
 wire \ann.bias[15] ;
 wire \ann.bias[16] ;
 wire \ann.bias[17] ;
 wire \ann.bias[18] ;
 wire \ann.bias[19] ;
 wire \ann.bias[1] ;
 wire \ann.bias[20] ;
 wire \ann.bias[21] ;
 wire \ann.bias[22] ;
 wire \ann.bias[23] ;
 wire \ann.bias[24] ;
 wire \ann.bias[25] ;
 wire \ann.bias[26] ;
 wire \ann.bias[27] ;
 wire \ann.bias[28] ;
 wire \ann.bias[29] ;
 wire \ann.bias[2] ;
 wire \ann.bias[30] ;
 wire \ann.bias[31] ;
 wire \ann.bias[3] ;
 wire \ann.bias[4] ;
 wire \ann.bias[5] ;
 wire \ann.bias[6] ;
 wire \ann.bias[7] ;
 wire \ann.bias[8] ;
 wire \ann.bias[9] ;
 wire \ann.in_ff[0][0] ;
 wire \ann.in_ff[0][10] ;
 wire \ann.in_ff[0][11] ;
 wire \ann.in_ff[0][12] ;
 wire \ann.in_ff[0][13] ;
 wire \ann.in_ff[0][14] ;
 wire \ann.in_ff[0][15] ;
 wire \ann.in_ff[0][1] ;
 wire \ann.in_ff[0][2] ;
 wire \ann.in_ff[0][3] ;
 wire \ann.in_ff[0][4] ;
 wire \ann.in_ff[0][5] ;
 wire \ann.in_ff[0][6] ;
 wire \ann.in_ff[0][7] ;
 wire \ann.in_ff[0][8] ;
 wire \ann.in_ff[0][9] ;
 wire \ann.in_ff[1][0] ;
 wire \ann.in_ff[1][10] ;
 wire \ann.in_ff[1][11] ;
 wire \ann.in_ff[1][12] ;
 wire \ann.in_ff[1][13] ;
 wire \ann.in_ff[1][14] ;
 wire \ann.in_ff[1][15] ;
 wire \ann.in_ff[1][1] ;
 wire \ann.in_ff[1][2] ;
 wire \ann.in_ff[1][3] ;
 wire \ann.in_ff[1][4] ;
 wire \ann.in_ff[1][5] ;
 wire \ann.in_ff[1][6] ;
 wire \ann.in_ff[1][7] ;
 wire \ann.in_ff[1][8] ;
 wire \ann.in_ff[1][9] ;
 wire \ann.in_ff[2][0] ;
 wire \ann.in_ff[2][10] ;
 wire \ann.in_ff[2][11] ;
 wire \ann.in_ff[2][12] ;
 wire \ann.in_ff[2][13] ;
 wire \ann.in_ff[2][14] ;
 wire \ann.in_ff[2][15] ;
 wire \ann.in_ff[2][1] ;
 wire \ann.in_ff[2][2] ;
 wire \ann.in_ff[2][3] ;
 wire \ann.in_ff[2][4] ;
 wire \ann.in_ff[2][5] ;
 wire \ann.in_ff[2][6] ;
 wire \ann.in_ff[2][7] ;
 wire \ann.in_ff[2][8] ;
 wire \ann.in_ff[2][9] ;
 wire \ann.ldX ;
 wire \ann.multiply_FF[0] ;
 wire \ann.multiply_FF[10] ;
 wire \ann.multiply_FF[11] ;
 wire \ann.multiply_FF[12] ;
 wire \ann.multiply_FF[13] ;
 wire \ann.multiply_FF[14] ;
 wire \ann.multiply_FF[15] ;
 wire \ann.multiply_FF[16] ;
 wire \ann.multiply_FF[17] ;
 wire \ann.multiply_FF[18] ;
 wire \ann.multiply_FF[19] ;
 wire \ann.multiply_FF[1] ;
 wire \ann.multiply_FF[20] ;
 wire \ann.multiply_FF[21] ;
 wire \ann.multiply_FF[22] ;
 wire \ann.multiply_FF[23] ;
 wire \ann.multiply_FF[24] ;
 wire \ann.multiply_FF[25] ;
 wire \ann.multiply_FF[26] ;
 wire \ann.multiply_FF[27] ;
 wire \ann.multiply_FF[28] ;
 wire \ann.multiply_FF[29] ;
 wire \ann.multiply_FF[2] ;
 wire \ann.multiply_FF[30] ;
 wire \ann.multiply_FF[31] ;
 wire \ann.multiply_FF[3] ;
 wire \ann.multiply_FF[4] ;
 wire \ann.multiply_FF[5] ;
 wire \ann.multiply_FF[6] ;
 wire \ann.multiply_FF[7] ;
 wire \ann.multiply_FF[8] ;
 wire \ann.multiply_FF[9] ;
 wire \ann.multiply_out[0] ;
 wire \ann.multiply_out[10] ;
 wire \ann.multiply_out[11] ;
 wire \ann.multiply_out[12] ;
 wire \ann.multiply_out[13] ;
 wire \ann.multiply_out[14] ;
 wire \ann.multiply_out[15] ;
 wire \ann.multiply_out[16] ;
 wire \ann.multiply_out[17] ;
 wire \ann.multiply_out[18] ;
 wire \ann.multiply_out[19] ;
 wire \ann.multiply_out[1] ;
 wire \ann.multiply_out[20] ;
 wire \ann.multiply_out[21] ;
 wire \ann.multiply_out[22] ;
 wire \ann.multiply_out[23] ;
 wire \ann.multiply_out[24] ;
 wire \ann.multiply_out[25] ;
 wire \ann.multiply_out[26] ;
 wire \ann.multiply_out[27] ;
 wire \ann.multiply_out[28] ;
 wire \ann.multiply_out[29] ;
 wire \ann.multiply_out[2] ;
 wire \ann.multiply_out[30] ;
 wire \ann.multiply_out[31] ;
 wire \ann.multiply_out[3] ;
 wire \ann.multiply_out[4] ;
 wire \ann.multiply_out[5] ;
 wire \ann.multiply_out[6] ;
 wire \ann.multiply_out[7] ;
 wire \ann.multiply_out[8] ;
 wire \ann.multiply_out[9] ;
 wire \ann.next_state[0] ;
 wire \ann.next_state[1] ;
 wire \ann.state[0] ;
 wire \ann.state[1] ;
 wire \ann.sum[0] ;
 wire \ann.sum[10] ;
 wire \ann.sum[11] ;
 wire \ann.sum[12] ;
 wire \ann.sum[13] ;
 wire \ann.sum[14] ;
 wire \ann.sum[15] ;
 wire \ann.sum[16] ;
 wire \ann.sum[17] ;
 wire \ann.sum[18] ;
 wire \ann.sum[19] ;
 wire \ann.sum[1] ;
 wire \ann.sum[20] ;
 wire \ann.sum[21] ;
 wire \ann.sum[22] ;
 wire \ann.sum[23] ;
 wire \ann.sum[24] ;
 wire \ann.sum[25] ;
 wire \ann.sum[26] ;
 wire \ann.sum[27] ;
 wire \ann.sum[28] ;
 wire \ann.sum[29] ;
 wire \ann.sum[2] ;
 wire \ann.sum[30] ;
 wire \ann.sum[31] ;
 wire \ann.sum[3] ;
 wire \ann.sum[4] ;
 wire \ann.sum[5] ;
 wire \ann.sum[6] ;
 wire \ann.sum[7] ;
 wire \ann.sum[8] ;
 wire \ann.sum[9] ;
 wire \ann.temp[0] ;
 wire \ann.temp[10] ;
 wire \ann.temp[11] ;
 wire \ann.temp[12] ;
 wire \ann.temp[13] ;
 wire \ann.temp[14] ;
 wire \ann.temp[15] ;
 wire \ann.temp[16] ;
 wire \ann.temp[17] ;
 wire \ann.temp[18] ;
 wire \ann.temp[19] ;
 wire \ann.temp[1] ;
 wire \ann.temp[20] ;
 wire \ann.temp[21] ;
 wire \ann.temp[22] ;
 wire \ann.temp[23] ;
 wire \ann.temp[24] ;
 wire \ann.temp[25] ;
 wire \ann.temp[26] ;
 wire \ann.temp[27] ;
 wire \ann.temp[28] ;
 wire \ann.temp[29] ;
 wire \ann.temp[2] ;
 wire \ann.temp[30] ;
 wire \ann.temp[3] ;
 wire \ann.temp[4] ;
 wire \ann.temp[5] ;
 wire \ann.temp[6] ;
 wire \ann.temp[7] ;
 wire \ann.temp[8] ;
 wire \ann.temp[9] ;
 wire \ann.weight[0] ;
 wire \ann.weight[10] ;
 wire \ann.weight[11] ;
 wire \ann.weight[12] ;
 wire \ann.weight[13] ;
 wire \ann.weight[14] ;
 wire \ann.weight[15] ;
 wire \ann.weight[1] ;
 wire \ann.weight[2] ;
 wire \ann.weight[3] ;
 wire \ann.weight[4] ;
 wire \ann.weight[5] ;
 wire \ann.weight[6] ;
 wire \ann.weight[7] ;
 wire \ann.weight[8] ;
 wire \ann.weight[9] ;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net22;
 wire net223;
 wire net23;
 wire net24;
 wire net25;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__A (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(\ann.temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A (.DIODE(\ann.ReLU_out[1][22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__D (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__D (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__C1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__C1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__C (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__D (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__C (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A2 (.DIODE(\ann.weight[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__C (.DIODE(\ann.weight[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B (.DIODE(\ann.weight[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__C1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A (.DIODE(\ann.in_ff[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__B2 (.DIODE(\ann.in_ff[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__B (.DIODE(\ann.in_ff[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__C1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__C (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__C (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A (.DIODE(\ann.in_ff[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__B (.DIODE(\ann.weight[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A2 (.DIODE(\ann.weight[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__C (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A1_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A2_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__C (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(\ann.in_ff[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A1 (.DIODE(\ann.in_ff[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A2 (.DIODE(\ann.weight[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B1 (.DIODE(\ann.weight[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B2 (.DIODE(\ann.in_ff[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__D (.DIODE(\ann.weight[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B (.DIODE(\ann.weight[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A2 (.DIODE(\ann.weight[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__D (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__C (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A1_N (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A2_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A1 (.DIODE(\ann.in_ff[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A (.DIODE(\ann.in_ff[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__C (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__D (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A1_N (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A2_N (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A (.DIODE(\ann.in_ff[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A2 (.DIODE(\ann.weight[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B1 (.DIODE(\ann.weight[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__D (.DIODE(\ann.weight[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__B (.DIODE(\ann.in_ff[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__D (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A2_N (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A (.DIODE(\ann.in_ff[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__C (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__D (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A2_N (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__C (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A1_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A2_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__C (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__C (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__D (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A1_N (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A2_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B (.DIODE(\ann.weight[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__D (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__C (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__D (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__D (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A2_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__B (.DIODE(\ann.weight[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__C (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__C1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__B1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__C (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__C (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__D (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__D (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A1_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A2_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__C (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B1 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__C (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__D (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__C (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__C (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__D (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1_N (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A_N (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__C (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__D (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__D (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__C (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__C (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__D (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__C (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__D (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__C (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__D (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__D (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1_N (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A2_N (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__C (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(\ann.weight[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__C (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__B1_N (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__C (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__D (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__C (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__D (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A2_N (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__D (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__C (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A1_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A2_N (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__B (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A_N (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__C (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__C (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A (.DIODE(_1918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A (.DIODE(_1918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__C (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(\ann.in_ff[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A (.DIODE(\ann.in_ff[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__C (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A2 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A (.DIODE(\ann.in_ff[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__C (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__C (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(\ann.in_ff[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A (.DIODE(\ann.in_ff[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__D (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__C (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A1 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A1 (.DIODE(\ann.in_ff[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A_N (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__B (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A_N (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__B (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__C (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__D (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__B (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B (.DIODE(_1918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__B (.DIODE(_1918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A (.DIODE(\ann.in_ff[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__C (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__C (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__B (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__B (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__B (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__B (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A1 (.DIODE(\ann.in_ff[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A3 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A4 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A2 (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__B1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__C (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A1_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A2_N (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__D (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A1 (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__B (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__C (.DIODE(\ann.weight[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__C (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A_N (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__B (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A2 (.DIODE(_2409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A1 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__B (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A_N (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A1 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A (.DIODE(_1918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A (.DIODE(_1918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__B (.DIODE(\ann.weight[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A_N (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__B (.DIODE(_2497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A1 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__B (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__C (.DIODE(\ann.weight[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__C (.DIODE(\ann.weight[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A_N (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A (.DIODE(_2222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A_N (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B (.DIODE(_2505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A (.DIODE(_2505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A (.DIODE(_1360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__B1 (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A1 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A_N (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A2 (.DIODE(\ann.weight[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__B (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__B (.DIODE(_2654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A1 (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A0 (.DIODE(_2226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A1 (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B (.DIODE(_2696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A1 (.DIODE(\ann.multiply_FF[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B (.DIODE(\ann.multiply_FF[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(\ann.multiply_FF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__B (.DIODE(\ann.multiply_FF[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__C (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__B (.DIODE(\ann.sum[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__B (.DIODE(\ann.sum[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__B (.DIODE(\ann.sum[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B (.DIODE(\ann.sum[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(\ann.sum[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__C1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A (.DIODE(\ann.bias[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A (.DIODE(\ann.bias[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__C (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A1 (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__B (.DIODE(_3104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__B2 (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A1 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__B2 (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A2_N (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A2 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__B2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A2_N (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B2 (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__B (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__B (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__B1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B2 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__B2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__B1 (.DIODE(_3133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A1 (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A2 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A2_N (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A1 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A2 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__B1 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A2 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__B1 (.DIODE(_0584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__B2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A1_N (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__A2_N (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__B1 (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A2 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__A1 (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A1 (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A2 (.DIODE(_3226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A2_N (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__A (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A1 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__B1 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A2 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__B1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__B2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A1_N (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__A2_N (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B1 (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A2 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A1 (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A (.DIODE(\ann.temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A1 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A2 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B1 (.DIODE(_0602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A2_N (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__B2 (.DIODE(_0602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__B2 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__A1 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__A1 (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A1_N (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__B2 (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A1 (.DIODE(_3305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A1 (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__B2 (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__B1 (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A (.DIODE(\ann.temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__B2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__A1 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__B2 (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__B2 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__A2_N (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__B1 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__B1 (.DIODE(_0609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__A2 (.DIODE(_0609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__B1 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__A2 (.DIODE(_0610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__A1 (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__B2 (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__A1 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__A (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__B2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__A1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__B1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__A1 (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__B2 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A1 (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__B2 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__A2_N (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__B1 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__A1 (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__B2 (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__A1 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__B2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__B1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__A1 (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__B2 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__A1_N (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__B2 (.DIODE(\ann.temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__B2 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__A (.DIODE(_3487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__B2 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__B2 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__B2 (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__A1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__B1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__A1 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__B2 (.DIODE(\ann.temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__A1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__B2 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__A2_N (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__A1 (.DIODE(\ann.temp[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__B1 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__B2 (.DIODE(\ann.temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__A1 (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__B2 (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__A1 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__A (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__A (.DIODE(\ann.temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__B2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__A1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__B1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__A1 (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__B2 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__B2 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__A2 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__B2 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__A2 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__B1 (.DIODE(\ann.temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__A1 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__B2 (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__A2 (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__B1 (.DIODE(\ann.temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__A1 (.DIODE(_3587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__A2 (.DIODE(\ann.temp[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__B1 (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__B (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__A1 (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A2_N (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__B2 (.DIODE(\ann.temp[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__B (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__B (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__A1 (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__B2 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__A1 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__A1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__B2 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__B1 (.DIODE(\ann.ReLU_out[1][22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__B2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__A1 (.DIODE(_0580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__B1 (.DIODE(\ann.temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__A1 (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__A1 (.DIODE(\ann.temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__B1_N (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__A2 (.DIODE(_3632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__B1_N (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7288__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7290__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__S (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__S (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__S (.DIODE(_3384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7300__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7302__S (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7303__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7304__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7307__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7308__S (.DIODE(_3384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7309__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7310__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7313__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7316__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7317__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7319__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7323__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7324__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7328__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7330__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7331__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7334__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7338__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7340__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7341__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7342__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7344__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7345__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7346__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7347__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7348__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7349__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7351__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7352__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7353__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7355__S (.DIODE(_3566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7357__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7358__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7359__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7360__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7361__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7362__S (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7363__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7364__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7366__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7368__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7372__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7373__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__A0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7375__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7377__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7378__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7383__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7384__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7385__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7386__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7387__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7389__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7394__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7405__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7406__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7408__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7409__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7413__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7415__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7419__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7424__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7427__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7429__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7433__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7434__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7436__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7437__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7439__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7444__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7446__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7447__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7449__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7450__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7450__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7451__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__B1_N (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7453__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7454__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7460__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7461__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7463__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7463__B1_N (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7467__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7468__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7472__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7476__A0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__7476__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7479__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7480__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7483__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7486__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7488__S (.DIODE(_3566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7491__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7492__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7493__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7497__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7498__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7499__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__A0 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7502__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7503__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7504__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7505__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7506__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7507__A0 (.DIODE(\ann.ReLU_out[1][22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7507__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7508__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7509__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7510__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7511__A0 (.DIODE(_3842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7511__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7512__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7513__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7514__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7515__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7516__A0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__7516__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7517__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7518__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7520__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7521__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7523__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7524__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7525__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7526__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7528__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7529__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7530__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__7531__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__7532__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7533__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7534__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7535__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7536__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7537__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__7539__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7540__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7541__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7542__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7543__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__7544__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7545__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7546__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7547__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7549__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7550__S (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7551__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7552__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7553__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7554__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__7555__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__7557__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7558__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7560__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7561__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7562__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7566__S (.DIODE(_3637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7567__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7568__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7572__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7573__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7575__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7577__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7578__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7579__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7580__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7581__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7582__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7583__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7584__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7585__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7586__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7587__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__7588__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__7589__S (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7590__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__7591__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__7592__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7594__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__7595__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7598__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7599__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__7599__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__7600__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__7600__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7605__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7606__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7607__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7607__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7608__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7610__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7613__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7613__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7615__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7615__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7617__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7617__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7618__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7619__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7619__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7620__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7620__B (.DIODE(\ann.sum[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7622__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7622__B (.DIODE(\ann.sum[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7623__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7623__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7625__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7625__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7627__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7627__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7628__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7629__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7629__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7632__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7636__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7637__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7637__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7638__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__7639__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7639__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7642__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7643__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7643__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7644__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7645__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7645__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7646__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7647__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7647__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7648__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7650__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7651__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7652__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7653__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7653__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7654__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7655__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7655__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7656__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7657__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7657__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7658__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7659__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7659__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7660__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7661__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7661__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7662__A_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7663__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7663__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7665__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7665__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7666__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7667__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7667__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7668__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7668__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7670__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7670__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7671__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7671__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7672__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7672__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7673__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7673__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7674__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7674__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7675__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7675__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7676__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7676__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7677__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7677__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7678__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7678__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7680__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7680__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7681__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7681__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7684__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7684__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7685__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7685__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7686__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7686__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7687__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7687__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7688__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7688__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7689__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7690__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7690__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__7691__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7691__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7692__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7692__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7693__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7693__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7694__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7694__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7695__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7695__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__7696__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__7696__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__7696__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7697__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7697__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7698__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7699__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7699__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7700__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7700__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7701__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7701__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7702__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7702__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7704__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7704__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7705__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7705__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7706__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7706__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7709__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7709__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7710__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7710__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7711__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7711__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7712__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7712__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7713__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7713__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7714__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7714__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7715__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7715__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7716__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7716__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7717__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7717__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7718__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7718__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7719__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7719__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7720__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7720__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7721__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7722__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7722__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__7723__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7723__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7724__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7724__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7725__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7725__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7726__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7726__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7729__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7729__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7730__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7731__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7731__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7732__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7732__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7733__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7733__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7734__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7734__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7736__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7736__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7737__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7737__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7738__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7738__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7740__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7740__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7741__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7741__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7742__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7742__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7743__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7743__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7744__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7744__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7745__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7745__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7746__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7746__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7747__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7747__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7748__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7748__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7749__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7749__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7750__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7750__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7751__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7751__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7752__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7752__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7753__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7754__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7754__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__7755__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7755__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7757__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7757__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7758__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7758__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7759__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7759__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__7760__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__7760__C_N (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__7761__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__7761__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__7761__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7764__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7764__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7766__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7766__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7767__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7767__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7768__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7768__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7769__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7769__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7770__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7770__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7771__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7771__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7772__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7772__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7773__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7773__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7774__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7774__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7776__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7776__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7777__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7777__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7778__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7778__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7780__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7780__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7781__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7781__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7782__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7782__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7784__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7784__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7785__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7785__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7786__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__7787__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7787__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7792__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7792__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__7793__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__7793__C (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__7794__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__7794__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7796__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7798__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7798__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7799__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7799__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7800__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7800__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7802__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7802__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7803__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7803__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7804__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7804__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7805__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7805__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7806__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7806__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7807__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7807__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7808__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7808__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7809__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7809__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7810__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7810__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7813__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7813__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7814__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7814__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7815__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7815__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7816__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7816__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7817__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7817__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7818__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7818__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7819__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__7820__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7820__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7821__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7821__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7822__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7822__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7823__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7823__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7824__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7824__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7825__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7825__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__7826__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__7826__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__7827__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7827__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7828__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7829__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7829__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7830__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7830__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7831__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7831__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7832__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7832__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7834__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7834__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7835__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7835__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7836__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7836__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7837__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7837__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7838__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7838__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7839__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7839__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7840__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7840__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7841__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7841__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7842__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7842__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7843__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7843__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7844__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7844__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7845__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7845__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7846__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7846__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7847__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7847__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7848__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7848__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7849__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7849__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7850__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7850__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7851__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7852__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7852__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7853__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7853__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7854__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7854__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7856__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7856__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7857__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7857__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__7858__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__7859__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7859__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7860__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7861__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7861__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7862__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7862__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7863__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7863__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7864__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7864__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7865__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7865__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7867__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7867__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7868__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7868__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7869__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7869__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7871__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7871__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7872__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7872__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7874__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7874__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7875__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7875__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7876__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7876__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7878__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7878__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7880__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7880__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7881__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7881__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7882__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7882__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7883__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7884__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7884__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__7885__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7885__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7886__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7886__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7887__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7887__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7889__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7889__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__7890__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__7890__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7892__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7892__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7895__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7895__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7896__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7896__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7897__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7897__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7898__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7898__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7899__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7899__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7901__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7901__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7903__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7903__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7906__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7906__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7907__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7907__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7908__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7908__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7909__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7909__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7910__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7910__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7912__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7912__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7914__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7914__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7916__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7919__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7919__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__7920__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7920__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7921__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7921__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7922__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7922__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__7923__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7925__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7927__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7929__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__7931__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7933__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7934__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__7935__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7939__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__A1 (.DIODE(\ann.sum[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__A1 (.DIODE(\ann.sum[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7945__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7947__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7949__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7951__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7953__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7955__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7959__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7961__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7963__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7965__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7967__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7969__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7971__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7973__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7975__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7977__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7979__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7981__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__7985__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__7985__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7987__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__7987__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7988__A1 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7988__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7989__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7990__A1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7990__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7991__A1 (.DIODE(_3928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7991__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7992__A1 (.DIODE(_3929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7992__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7993__A1 (.DIODE(_3930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7993__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7994__A1 (.DIODE(_3931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7994__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__A1 (.DIODE(_3932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__7996__A1 (.DIODE(_3933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7996__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__A1 (.DIODE(_3934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__A1 (.DIODE(_3935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__A1 (.DIODE(_3936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__A1 (.DIODE(_3937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8001__A1 (.DIODE(_3938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8001__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8002__A1 (.DIODE(_3939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8002__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8003__A1 (.DIODE(_3940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8003__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__A1 (.DIODE(_3941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__A1 (.DIODE(_3942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__A1 (.DIODE(_3943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8007__A1 (.DIODE(_3944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8007__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__A1 (.DIODE(_3945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8009__A1 (.DIODE(_3946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8009__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__A1 (.DIODE(_3947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__A1 (.DIODE(_3948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__8012__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__8013__A1 (.DIODE(_3950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8013__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__8014__A1 (.DIODE(_3951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8014__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__8015__A1 (.DIODE(_3952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8015__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__8016__A1 (.DIODE(_3953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8016__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8017__A1 (.DIODE(_3954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8017__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8018__A1 (.DIODE(_3955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8018__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__8019__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__8019__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8020__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8021__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__8021__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8022__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8024__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8025__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__8025__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8026__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8027__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__8027__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8028__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8029__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__8029__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8030__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8031__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__8031__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8032__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8033__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__8033__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8034__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8035__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__8035__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8036__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8037__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__8037__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8038__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8039__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__8039__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8040__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8041__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__8041__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8043__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__8043__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8044__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8045__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__8045__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8047__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__8047__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8049__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__8049__S (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__8051__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__8051__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8052__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8054__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8055__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__8055__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8056__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8057__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__8057__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8058__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8059__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__8059__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8060__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8061__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__8061__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8062__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8063__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__8063__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8064__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__8065__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__8065__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8066__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__8067__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__8067__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8068__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8069__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__8069__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8070__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8071__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__8071__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8072__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8073__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__8073__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8074__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8075__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__8075__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8076__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8077__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__8077__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8081__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__8081__S (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__8083__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__8083__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8084__A_N (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__8086__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__8086__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8087__A_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__8089__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__8089__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8090__A_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8093__A_N (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__8095__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__8095__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8096__A_N (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__8096__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8097__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8098__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__8098__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8099__A_N (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__8099__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8100__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8101__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__8101__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8102__A_N (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__8102__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8103__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8104__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__8104__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__A_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8106__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8107__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__8107__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8108__A_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__8108__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8109__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8110__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__8110__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8111__A_N (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__8111__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8112__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8113__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__8113__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__A_N (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8115__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8117__A_N (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__8120__A_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__8120__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__8121__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__8122__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__8122__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8123__A_N (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__8125__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__8125__S (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8126__A_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__8127__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8128__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__8128__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__A_N (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8130__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__8131__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8132__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__8134__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8136__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8138__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8156__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8166__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__8166__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8168__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__8168__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8172__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__8174__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__8176__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__8178__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__8180__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__8182__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__8184__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__8186__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__8188__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__8188__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8190__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__8192__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__8194__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__8194__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__8196__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__8197__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8198__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8199__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8200__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8201__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8202__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8203__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8204__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8205__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8206__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8208__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8209__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8210__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8211__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8212__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8213__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8214__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8215__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8216__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8217__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8218__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8219__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8221__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8222__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8223__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8224__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8225__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8226__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8227__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8228__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8229__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8230__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8231__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8232__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8232__D (.DIODE(_0101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__D (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__D (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8235__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8236__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8237__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8238__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8239__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8240__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8241__GATE_N (.DIODE(_0066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8242__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8243__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8244__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8245__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8246__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8247__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8248__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8249__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8250__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8251__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8252__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8253__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8254__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8255__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8256__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8257__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8258__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8259__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8260__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8261__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8262__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8263__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8264__GATE_N (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__8265__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8266__GATE_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__8267__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8268__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8269__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8270__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8271__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8272__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8273__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8274__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8275__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8276__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8277__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8278__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8279__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8280__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8281__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8282__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8283__D (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8283__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8284__D (.DIODE(_0008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8284__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8285__GATE_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__8286__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8287__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8288__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8289__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8290__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8291__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8292__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8293__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8294__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8295__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8296__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8297__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8298__GATE_N (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__8299__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8300__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8301__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8302__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8303__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8304__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8305__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8306__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8307__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8308__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8309__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8310__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8311__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8314__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8315__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8316__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8317__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8318__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8319__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8320__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8321__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8322__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8323__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8324__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8325__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8326__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8327__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8330__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8331__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8332__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8333__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8334__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8335__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8336__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8337__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8338__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8339__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8340__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8341__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8342__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8344__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8345__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8346__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8347__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8348__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8349__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8350__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8351__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8352__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8353__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8354__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8355__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8356__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8357__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8358__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8359__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8360__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8362__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8363__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8364__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8365__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8367__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8368__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8369__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8370__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8371__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8372__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8373__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8374__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8375__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8376__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8377__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8378__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8379__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8380__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8381__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8382__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8383__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8384__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8385__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8387__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8388__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8389__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8390__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8391__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8392__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8393__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8394__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8395__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8396__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8397__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8398__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8399__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8400__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8401__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8402__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8403__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8404__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8405__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8406__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8407__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8408__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8409__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8410__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8411__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8412__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8413__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8414__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8415__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8416__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8417__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8418__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8419__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8420__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8422__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8423__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8424__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8425__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8426__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8427__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8428__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8429__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8430__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8431__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8432__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8433__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8434__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8435__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8436__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8437__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8438__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8439__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8440__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8441__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8442__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8443__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8444__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8445__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8446__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8447__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8448__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8449__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8450__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8451__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8452__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8453__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8454__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8455__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8456__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8457__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8458__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8459__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8460__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8462__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8463__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8464__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8465__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8466__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8467__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8468__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8469__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8470__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8471__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8472__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8473__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8474__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8475__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8476__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8477__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8478__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8479__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8480__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8481__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8482__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8483__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8484__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8485__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8486__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8487__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8488__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8489__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8490__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8491__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8492__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8493__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8494__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8495__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8496__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8497__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8498__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8499__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8500__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8501__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8502__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8503__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8504__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8505__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8506__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8507__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8508__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8509__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8510__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8511__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8512__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8513__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8516__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8518__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8519__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8520__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8521__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8522__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8523__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8524__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8525__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8526__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8527__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8528__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8529__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8530__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8531__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8532__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8533__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8534__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8535__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8536__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8537__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8538__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8541__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8542__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8543__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8544__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8545__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8549__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8550__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8551__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8552__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8553__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8554__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8555__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8557__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8558__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8560__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8561__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8562__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8563__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8564__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8565__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8566__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8567__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8568__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8569__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8570__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8571__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8572__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8573__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8574__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8575__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8576__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8580__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8581__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8582__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8583__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8584__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8585__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8586__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8587__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8588__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8589__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8590__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8591__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8592__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8593__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8594__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8595__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8596__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8598__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8599__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8600__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8601__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8602__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8603__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8604__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8605__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8606__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8607__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8608__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8609__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8611__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8612__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8613__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8614__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8615__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8616__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8617__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8618__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8619__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8621__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8622__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8623__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8624__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8625__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8626__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8627__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8628__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8629__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8630__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8631__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8632__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8633__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8634__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8635__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8636__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8637__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8638__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8639__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8640__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8641__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8642__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8643__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8644__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8645__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8646__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8647__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8648__CLK (.DIODE(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8649__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8650__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8651__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8652__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8653__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8654__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8655__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8656__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8657__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8659__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8660__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8661__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8662__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8663__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8664__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8665__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8666__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8667__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8668__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8669__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8670__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8671__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8672__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8674__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8675__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8676__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8677__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8678__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8679__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8680__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8681__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8682__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8683__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8684__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8685__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8686__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8687__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8688__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8689__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8690__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8691__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8692__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8693__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8694__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8695__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8696__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8697__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8698__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8699__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8700__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8701__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8702__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8703__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8704__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8705__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8706__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8706__D (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__8707__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8707__D (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__8708__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8708__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__8709__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8709__D (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__8710__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8710__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__8711__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8711__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__8712__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8712__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__8713__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8713__D (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__8714__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8714__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__8715__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8715__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__8716__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8716__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__8717__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8717__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__8719__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8719__D (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__8720__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8720__D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__D (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__8722__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8723__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8724__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8725__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8726__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8727__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8728__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8729__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8730__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8731__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8732__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8733__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8734__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8735__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8736__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8737__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8738__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8739__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8740__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8741__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8742__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8743__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8744__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8745__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8746__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8747__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8748__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8749__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8750__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8751__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8752__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8753__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8754__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8755__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8756__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8757__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8758__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8759__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8760__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8761__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8762__CLK (.DIODE(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8763__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8764__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8765__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8766__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8767__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8768__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8769__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(\ann.in_ff[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(\ann.weight[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(\ann.weight[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(\ann.weight[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(\ann.weight[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(\ann.weight[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(\ann.weight[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(\ann.weight[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(\ann.weight[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(\ann.weight[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(\ann.weight[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(_3566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(_3384_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(_0066_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_3637_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold330_A (.DIODE(\ann.in_ff[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold365_A (.DIODE(\ann.in_ff[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold376_A (.DIODE(\ann.in_ff[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold388_A (.DIODE(\ann.in_ff[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold407_A (.DIODE(\ann.in_ff[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold408_A (.DIODE(\ann.in_ff[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold458_A (.DIODE(\ann.temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold463_A (.DIODE(\ann.temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold489_A (.DIODE(\ann.temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold494_A (.DIODE(\ann.ReLU_out[1][22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold499_A (.DIODE(\ann.temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold501_A (.DIODE(\ann.temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold503_A (.DIODE(\ann.temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold504_A (.DIODE(\ann.temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold511_A (.DIODE(\ann.temp[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold520_A (.DIODE(\ann.temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold528_A (.DIODE(\ann.temp[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold530_A (.DIODE(\ann.temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold531_A (.DIODE(\ann.temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold533_A (.DIODE(\ann.bias[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold534_A (.DIODE(\ann.temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1000_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1000_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1000_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1000_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1000_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1000_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1000_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1000_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1000_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1000_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1000_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1000_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1000_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1000_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1000_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1001_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1001_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1001_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1001_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1001_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1001_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1001_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1001_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1001_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1001_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1002_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1002_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1002_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1002_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1002_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1002_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1002_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1002_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1003_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1003_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1003_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1003_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1003_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1003_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1003_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1003_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1003_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1003_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1003_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1003_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1003_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1003_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1003_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1003_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1004_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1004_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1004_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1004_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1004_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1004_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1004_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1004_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1004_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1004_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1004_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1004_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1004_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1004_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1004_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1005_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1005_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1005_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1005_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1005_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1005_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1005_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1005_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1005_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1005_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1006_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1006_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1006_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1006_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1006_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1006_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1006_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1006_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1006_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1006_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1006_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1006_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1006_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1006_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1006_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1007_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1007_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1007_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1007_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1007_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1007_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1007_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1007_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1007_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1008_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1008_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1008_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1008_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1008_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1008_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1008_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1008_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1008_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1008_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1008_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1008_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1008_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1008_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1008_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1009_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1010_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1010_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1010_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1010_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1010_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1010_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1010_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1010_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1010_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1010_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1010_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1010_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1010_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1010_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1010_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1011_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1011_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1011_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1011_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1011_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1011_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1011_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1011_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1011_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1011_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1011_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1011_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1011_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1011_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1011_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1012_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1012_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1012_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1012_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1012_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1012_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1012_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1012_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1012_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1012_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1012_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1012_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1012_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1012_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1012_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1013_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1013_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1013_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1013_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1013_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1013_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1013_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1013_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1013_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1013_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1014_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1014_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1014_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1014_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1014_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1014_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1014_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1014_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1014_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1014_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1014_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1014_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1014_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1014_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1014_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1015_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1015_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1015_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1015_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1015_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1015_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1015_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1015_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1015_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1016_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1016_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1016_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1016_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1016_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1016_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1016_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1016_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1017_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1017_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1017_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1017_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1017_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1017_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1017_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1017_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1017_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1017_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1017_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1017_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1017_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1017_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1017_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1017_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1018_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1018_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1018_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1018_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1018_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1018_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1018_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1018_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1018_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1018_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1018_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1018_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1018_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1018_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1018_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1019_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1019_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1019_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1019_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1019_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1019_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1019_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1019_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1019_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1020_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1020_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1020_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1020_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1020_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1020_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1020_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1020_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1020_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1020_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1020_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1020_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1020_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1020_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1021_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1021_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1021_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1021_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1021_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1021_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1021_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1021_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1021_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1021_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1021_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1021_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1021_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1021_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1021_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1022_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1022_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1022_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1022_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1022_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1022_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1022_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1022_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1022_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1022_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1022_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1022_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1022_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1022_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1022_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1023_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1023_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1023_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1023_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1023_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1023_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1023_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1023_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1023_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1023_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1023_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1023_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1023_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1023_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1023_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1023_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1024_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1024_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1024_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1024_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1024_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1024_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1024_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1024_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1024_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1024_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1024_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1024_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1024_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1024_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1024_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1025_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1025_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1025_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1025_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1025_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1025_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1025_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1025_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1025_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1025_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1026_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1026_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1026_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1026_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1026_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1026_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1026_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1026_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1026_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1027_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1027_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1027_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1027_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1027_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1027_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1027_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1027_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1027_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1027_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1027_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1027_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1027_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1027_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1027_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1027_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1028_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1028_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1028_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1028_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1028_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1028_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1028_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1028_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1028_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1028_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1028_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1028_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1028_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1028_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1028_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1029_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1029_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1029_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1029_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1029_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1029_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1029_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1029_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1029_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1030_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1030_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1030_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1030_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1030_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1030_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1030_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1030_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1030_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1031_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1031_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1031_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1031_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1031_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1031_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1031_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1031_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1031_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1031_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1032_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1032_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1032_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1032_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1032_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1032_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1032_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1032_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1032_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1032_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1032_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1032_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1032_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1032_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1032_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1033_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1033_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1033_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1033_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1033_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1033_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1033_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1033_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1033_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1034_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1034_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1034_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1034_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1034_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1034_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1034_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1034_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1034_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1034_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1034_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1034_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1034_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1034_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1034_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1035_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1035_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1035_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1035_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1035_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1035_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1035_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1035_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1035_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1036_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1036_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1036_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1036_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1036_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1036_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1036_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1036_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1036_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1036_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1036_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1036_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1036_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1036_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1036_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1037_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1037_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1037_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1037_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1037_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1037_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1037_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1037_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1038_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1038_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1038_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1038_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1038_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1038_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1038_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1038_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1038_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1038_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1038_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1038_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1038_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1038_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1038_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1039_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1039_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1039_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1039_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1039_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1039_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1039_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1039_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1039_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1039_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1039_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1039_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1039_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1039_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1039_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1039_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1040_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1040_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1040_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1040_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1040_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1040_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1040_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1040_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1040_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1040_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1040_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1040_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1040_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1040_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1040_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1041_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1041_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1041_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1041_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1041_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1041_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1041_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1041_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1041_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1041_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1042_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1042_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1042_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1042_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1042_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1042_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1042_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1042_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1042_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1042_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1042_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1042_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1042_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1042_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1043_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1043_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1043_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1043_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1043_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1043_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1043_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1043_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1043_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1043_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1043_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1043_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1043_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1043_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1043_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1044_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1044_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1044_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1044_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1044_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1044_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1044_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1044_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1044_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1045_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1045_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1045_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1045_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1045_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1045_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1045_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1045_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1045_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1046_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1046_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1046_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1046_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1046_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1046_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1046_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1046_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1046_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1046_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1046_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1046_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1046_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1046_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1046_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1047_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1047_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1047_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1047_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1047_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1047_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1047_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1047_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1047_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1047_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1047_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1047_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1047_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1047_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1047_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1048_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1048_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1048_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1048_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1048_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1048_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1048_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1048_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1048_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1048_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1048_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1048_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1048_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1048_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1048_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1049_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1049_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1049_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1049_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1049_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1049_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1049_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1049_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1050_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1050_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1050_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1050_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1050_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1050_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1050_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1050_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1050_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1050_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1051_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1051_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1051_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1051_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1051_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1051_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1051_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1051_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1051_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1051_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1051_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1051_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1051_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1051_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1051_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1052_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1052_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1052_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1052_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1052_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1052_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1052_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1052_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1052_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1052_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1052_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1052_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1052_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1052_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1053_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1053_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1053_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1053_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1053_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1053_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1053_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1053_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1053_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1053_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1054_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1054_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1054_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1054_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1054_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1054_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1054_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1054_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1054_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1055_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1055_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1055_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1055_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1055_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1055_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1055_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1055_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1055_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1055_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1056_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1056_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1056_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1056_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1056_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1056_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1056_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1056_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1056_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1056_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1056_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1056_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1056_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1056_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1056_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1057_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1057_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1057_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1057_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1057_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1057_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1057_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1057_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1057_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1057_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1057_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1057_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1057_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1057_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1057_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1057_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1058_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1058_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1059_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1059_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1059_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1059_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1059_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1059_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1059_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1059_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1059_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1059_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1059_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1059_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1059_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1059_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1059_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1059_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1060_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1060_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1060_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1060_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1060_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1060_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1060_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1060_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1060_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1061_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1061_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1061_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1061_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1061_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1061_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1061_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1061_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1061_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1061_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1061_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1061_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1061_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1061_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1061_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1061_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1062_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1062_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1062_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1062_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1062_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1062_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1062_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1062_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1062_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1062_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1062_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1062_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1062_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1062_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1062_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1063_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1063_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1063_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1063_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1063_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1063_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1063_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1063_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1063_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1064_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1064_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1064_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1064_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1064_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1064_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1064_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1064_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1064_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1064_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1064_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1064_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1064_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1064_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1064_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1065_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1065_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1065_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1065_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1065_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1065_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1065_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1065_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1066_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1066_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1066_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1066_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1066_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1066_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1066_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1066_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1066_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1066_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1066_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1066_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1066_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1066_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1066_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1067_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1067_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1067_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1067_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1067_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1067_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1067_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1067_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1067_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1067_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1067_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1067_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1067_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1067_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1067_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1067_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1068_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1068_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1068_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1068_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1068_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1068_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1068_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1068_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1068_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1068_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1068_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1068_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1068_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1068_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1068_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1069_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1069_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1069_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1069_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1069_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1069_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1069_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1069_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1069_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1069_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1069_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1069_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1069_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1069_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1069_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1069_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1070_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1070_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1070_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1070_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1070_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1070_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1070_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1070_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1070_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1070_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1070_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1070_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1070_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1070_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1070_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1071_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1071_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1071_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1071_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1071_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1071_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1071_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1071_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1071_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1072_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1072_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1072_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1072_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1072_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1072_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1072_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1072_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1072_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1072_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1072_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1072_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1072_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1072_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1072_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1073_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1073_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1073_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1073_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1073_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1073_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1073_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1073_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1073_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1073_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1073_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1073_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1073_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1073_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1073_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1074_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1074_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1074_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1074_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1074_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1074_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1074_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1074_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1074_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1074_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1074_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1074_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1074_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1074_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1074_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1075_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1075_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1075_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1075_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1075_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1075_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1075_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1075_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1075_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1075_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1075_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1075_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1075_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1075_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1075_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1076_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1076_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1076_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1076_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1076_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1076_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1076_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1076_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1076_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1076_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1076_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1076_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1076_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1076_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1076_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1077_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1077_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1077_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1077_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1077_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1077_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1077_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1077_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1077_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1077_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1077_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1077_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1077_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1077_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1077_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1078_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1078_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1078_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1078_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1078_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1078_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1078_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1078_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1078_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1078_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1078_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1078_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1078_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1078_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1078_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1079_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1079_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1079_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1079_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1079_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1079_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1079_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1079_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1079_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1080_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1080_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1080_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1081_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1081_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1081_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1081_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1081_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1081_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1081_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1081_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1081_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1081_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1081_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1082_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1082_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1082_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1082_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1082_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1082_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1082_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1082_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1082_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1082_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1082_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1082_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1082_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1082_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1082_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1083_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1083_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1083_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1083_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1083_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1083_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1083_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1083_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1083_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1083_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1083_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1083_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1083_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1083_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1083_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1083_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1084_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1084_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1084_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1084_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1084_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1084_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1084_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1084_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1084_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1084_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1084_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1084_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1084_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1084_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1084_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1085_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1085_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1085_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1086_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1086_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1086_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1086_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1086_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1086_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1086_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1086_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1087_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1087_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1087_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1087_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1087_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1087_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1087_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1087_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1087_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1087_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1087_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1087_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1087_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1087_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1087_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1087_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1088_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1088_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1088_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1088_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1088_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1088_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1088_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1088_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1088_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1088_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1088_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1088_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1088_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1088_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1088_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1089_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1089_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1089_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1089_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1089_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1089_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1089_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1089_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1089_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1089_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1089_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1089_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1089_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1089_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1089_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1089_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1090_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1090_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1090_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1090_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1090_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1090_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1090_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1090_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1090_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1090_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1090_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1090_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1090_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1090_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1090_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1091_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1091_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1091_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1091_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1091_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1091_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1091_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1091_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1091_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1092_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1092_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1092_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1092_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1092_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1092_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1092_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1092_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1092_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1092_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1092_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1092_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1092_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1092_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1092_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1093_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_251_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_269_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_279_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_283_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_287_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_288_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_291_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_293_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_295_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_297_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_299_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_301_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_301_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_303_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_305_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_305_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_307_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_307_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_307_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_311_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_311_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_313_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_315_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_317_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_317_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_319_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_323_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_325_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_327_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_327_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_329_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_329_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_331_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_333_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_333_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_335_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_335_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_337_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_339_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_339_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_341_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_343_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_345_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_345_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_347_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_349_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_351_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_353_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_355_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_357_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_357_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_358_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_359_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_359_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_359_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_359_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_359_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_360_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_360_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_360_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_361_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_361_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_361_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_361_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_362_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_362_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_362_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_363_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_363_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_363_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_363_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_364_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_364_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_364_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_366_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_366_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_366_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_367_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_367_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_367_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_367_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_368_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_368_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_368_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_369_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_370_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_370_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_370_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_371_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_371_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_371_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_372_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_372_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_372_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_373_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_373_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_373_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_374_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_374_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_375_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_375_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_376_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_377_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_377_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_378_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_379_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_379_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_380_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_380_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_380_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_381_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_381_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_381_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_381_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_382_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_382_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_382_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_383_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_383_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_383_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_383_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_383_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_384_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_384_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_385_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_385_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_385_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_386_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_387_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_387_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_387_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_387_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_388_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_388_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_388_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_389_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_389_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_389_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_389_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_390_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_390_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_390_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_391_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_391_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_391_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_391_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_392_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_392_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_392_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_392_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_392_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_392_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_394_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_394_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_394_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_394_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_394_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_394_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_395_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_395_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_395_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_395_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_395_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_395_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_395_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_395_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_395_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_395_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_395_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_395_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_395_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_396_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_396_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_396_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_396_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_396_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_396_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_396_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_396_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_397_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_397_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_397_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_397_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_397_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_397_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_397_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_397_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_398_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_398_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_398_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_398_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_398_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_398_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_398_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_398_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_398_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_398_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_398_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_399_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_399_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_399_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_399_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_399_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_399_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_399_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_399_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_399_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_400_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_400_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_400_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_400_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_400_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_400_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_401_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_401_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_401_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_401_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_401_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_401_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_401_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_402_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_402_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_402_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_402_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_402_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_402_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_402_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_402_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_402_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_402_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_402_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_402_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_402_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_402_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_402_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_402_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_402_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_402_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_403_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_403_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_403_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_403_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_403_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_403_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_403_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_403_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_403_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_403_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_403_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_403_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_404_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_404_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_404_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_404_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_404_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_404_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_404_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_404_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_404_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_404_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_405_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_405_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_405_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_405_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_405_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_405_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_405_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_406_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_406_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_406_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_406_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_407_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_407_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_407_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_407_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_407_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_407_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_407_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_408_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_408_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_408_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_408_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_408_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_408_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_408_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_408_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_408_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_408_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_408_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_408_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_408_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_409_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_409_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_409_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_409_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_409_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_409_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_409_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_409_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_409_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_409_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_409_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_409_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_409_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_410_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_410_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_410_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_410_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_410_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_410_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_410_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_410_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_410_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_410_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_411_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_411_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_411_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_411_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_411_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_411_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_411_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_411_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_411_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_411_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_412_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_412_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_412_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_412_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_412_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_412_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_412_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_412_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_412_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_413_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_413_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_413_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_413_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_413_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_413_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_413_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_413_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_413_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_413_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_413_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_414_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_414_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_414_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_414_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_414_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_414_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_414_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_414_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_414_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_415_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_415_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_415_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_415_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_415_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_415_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_415_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_415_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_415_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_416_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_416_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_416_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_416_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_416_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_416_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_416_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_416_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_416_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_416_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_416_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_416_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_416_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_416_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_416_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_416_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_417_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_417_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_417_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_417_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_417_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_417_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_417_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_417_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_417_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_418_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_418_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_418_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_418_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_418_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_418_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_418_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_418_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_418_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_418_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_418_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_418_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_418_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_419_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_419_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_419_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_419_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_419_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_419_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_419_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_419_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_419_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_419_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_420_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_420_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_420_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_420_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_420_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_420_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_420_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_420_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_420_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_420_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_420_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_420_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_421_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_421_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_421_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_421_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_421_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_421_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_421_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_422_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_422_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_422_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_422_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_422_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_422_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_422_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_422_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_422_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_423_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_423_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_423_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_423_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_423_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_423_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_423_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_423_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_423_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_423_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_423_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_423_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_423_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_423_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_423_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_423_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_424_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_424_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_424_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_424_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_424_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_424_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_424_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_424_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_424_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_424_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_424_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_424_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_425_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_425_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_425_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_425_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_425_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_425_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_425_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_425_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_425_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_425_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_425_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_425_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_426_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_426_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_426_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_426_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_426_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_426_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_426_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_426_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_426_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_426_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_426_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_426_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_426_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_426_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_427_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_427_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_427_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_427_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_427_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_427_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_427_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_427_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_427_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_427_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_427_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_427_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_427_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_428_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_428_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_428_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_428_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_428_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_428_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_428_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_428_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_428_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_428_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_428_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_428_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_428_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_428_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_428_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_429_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_429_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_429_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_429_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_429_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_429_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_429_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_429_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_429_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_429_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_429_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_430_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_430_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_430_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_430_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_430_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_430_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_430_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_430_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_430_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_430_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_430_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_430_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_430_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_431_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_431_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_431_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_431_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_431_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_431_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_431_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_431_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_431_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_431_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_431_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_431_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_432_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_432_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_432_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_432_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_432_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_432_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_432_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_432_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_432_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_432_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_432_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_432_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_433_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_433_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_433_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_433_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_433_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_433_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_434_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_434_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_434_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_434_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_434_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_434_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_434_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_435_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_435_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_435_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_435_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_435_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_435_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_435_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_435_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_435_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_436_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_436_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_436_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_436_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_436_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_436_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_436_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_436_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_436_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_436_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_436_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_436_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_436_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_436_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_436_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_437_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_437_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_437_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_437_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_437_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_437_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_437_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_437_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_437_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_437_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_437_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_437_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_438_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_438_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_438_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_438_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_439_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_439_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_439_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_439_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_439_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_439_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_439_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_439_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_440_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_440_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_440_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_440_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_440_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_440_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_440_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_440_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_441_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_441_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_441_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_441_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_441_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_441_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_441_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_441_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_441_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_441_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_441_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_441_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_441_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_441_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_441_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_442_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_442_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_442_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_442_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_442_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_442_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_442_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_442_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_442_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_442_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_442_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_442_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_442_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_442_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_442_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_442_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_442_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_442_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_442_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_443_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_443_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_443_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_443_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_443_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_443_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_443_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_443_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_443_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_443_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_443_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_443_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_443_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_444_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_444_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_444_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_444_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_444_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_444_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_444_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_444_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_444_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_444_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_444_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_444_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_444_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_444_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_444_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_444_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_444_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_444_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_445_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_445_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_445_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_445_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_445_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_445_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_445_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_445_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_445_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_445_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_445_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_445_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_446_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_446_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_446_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_446_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_446_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_446_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_447_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_447_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_447_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_447_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_447_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_448_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_448_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_448_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_448_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_448_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_448_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_449_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_449_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_449_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_450_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_450_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_450_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_450_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_450_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_450_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_450_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_450_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_450_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_450_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_450_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_450_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_450_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_450_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_450_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_450_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_450_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_450_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_450_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_451_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_451_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_451_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_451_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_451_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_451_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_451_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_451_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_451_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_451_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_451_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_451_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_451_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_451_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_451_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_452_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_452_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_452_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_452_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_452_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_452_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_452_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_452_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_452_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_452_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_452_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_452_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_453_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_453_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_453_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_453_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_453_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_453_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_453_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_453_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_453_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_453_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_453_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_454_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_454_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_454_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_454_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_455_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_455_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_455_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_455_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_455_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_455_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_455_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_456_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_456_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_456_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_456_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_456_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_456_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_457_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_457_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_457_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_457_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_457_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_457_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_457_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_457_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_457_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_457_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_458_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_458_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_458_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_458_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_458_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_458_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_458_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_458_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_458_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_459_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_459_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_459_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_459_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_459_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_459_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_459_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_459_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_460_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_460_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_460_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_460_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_460_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_460_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_460_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_460_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_460_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_460_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_460_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_460_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_460_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_460_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_460_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_460_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_461_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_461_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_461_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_461_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_461_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_461_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_461_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_462_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_462_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_462_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_462_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_462_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_462_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_462_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_462_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_462_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_462_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_462_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_462_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_462_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_462_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_462_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_462_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_462_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_463_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_463_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_463_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_463_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_463_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_463_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_463_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_463_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_463_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_463_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_463_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_463_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_464_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_464_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_464_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_464_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_464_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_464_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_464_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_464_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_464_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_464_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_464_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_464_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_464_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_464_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_464_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_465_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_465_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_465_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_465_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_465_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_465_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_466_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_466_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_466_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_466_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_466_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_466_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_466_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_466_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_466_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_466_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_467_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_467_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_467_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_467_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_467_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_467_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_467_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_468_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_468_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_468_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_468_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_468_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_468_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_468_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_468_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_468_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_468_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_468_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_468_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_468_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_468_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_468_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_469_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_469_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_469_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_469_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_469_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_469_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_469_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_469_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_469_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_469_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_469_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_469_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_469_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_469_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_469_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_469_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_470_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_470_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_470_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_470_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_470_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_470_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_470_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_470_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_470_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_470_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_470_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_470_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_471_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_471_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_471_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_471_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_471_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_471_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_471_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_471_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_472_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_472_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_472_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_472_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_472_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_472_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_472_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_472_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_472_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_472_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_472_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_472_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_472_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_472_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_473_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_473_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_473_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_473_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_473_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_473_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_473_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_473_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_473_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_474_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_474_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_474_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_474_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_474_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_474_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_474_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_474_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_474_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_474_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_474_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_475_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_475_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_475_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_475_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_475_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_475_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_475_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_476_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_476_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_476_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_476_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_476_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_476_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_477_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_477_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_478_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_478_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_478_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_478_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_478_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_478_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_478_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_478_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_478_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_478_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_479_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_479_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_479_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_479_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_479_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_479_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_479_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_479_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_480_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_480_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_480_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_480_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_480_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_480_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_480_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_480_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_480_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_480_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_480_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_480_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_481_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_481_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_481_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_481_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_481_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_481_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_481_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_481_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_481_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_482_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_482_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_482_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_482_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_482_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_482_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_482_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_482_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_483_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_483_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_483_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_483_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_483_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_483_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_483_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_483_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_483_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_484_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_484_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_484_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_484_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_484_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_484_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_484_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_484_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_484_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_484_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_484_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_484_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_484_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_484_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_484_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_484_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_484_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_485_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_485_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_485_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_485_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_485_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_485_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_485_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_486_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_486_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_486_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_486_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_486_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_486_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_486_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_486_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_486_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_486_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_486_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_486_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_486_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_486_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_487_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_487_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_487_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_487_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_487_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_487_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_487_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_487_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_487_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_487_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_487_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_487_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_487_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_487_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_488_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_488_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_488_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_488_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_488_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_488_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_488_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_488_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_488_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_488_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_489_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_489_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_489_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_489_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_489_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_489_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_489_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_489_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_489_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_489_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_489_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_489_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_490_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_490_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_490_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_490_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_490_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_490_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_490_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_490_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_490_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_490_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_490_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_490_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_491_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_491_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_491_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_491_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_491_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_491_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_492_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_492_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_492_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_492_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_492_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_492_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_492_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_492_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_493_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_493_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_493_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_493_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_493_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_493_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_493_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_493_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_493_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_493_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_493_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_493_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_493_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_493_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_493_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_494_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_494_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_494_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_494_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_494_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_494_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_494_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_494_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_494_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_494_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_494_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_494_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_494_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_494_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_494_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_495_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_495_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_495_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_495_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_495_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_495_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_496_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_496_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_496_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_496_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_496_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_496_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_496_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_496_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_496_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_496_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_496_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_496_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_496_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_497_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_497_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_497_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_497_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_497_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_498_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_498_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_498_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_498_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_498_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_498_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_498_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_498_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_498_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_498_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_498_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_498_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_498_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_498_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_498_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_498_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_498_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_498_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_498_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_498_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_498_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_498_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_498_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_499_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_499_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_499_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_499_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_499_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_499_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_499_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_499_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_500_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_500_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_500_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_500_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_500_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_500_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_500_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_500_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_500_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_500_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_500_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_500_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_500_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_500_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_500_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_500_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_500_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_500_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_500_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_500_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_500_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_500_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_501_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_501_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_501_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_501_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_501_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_501_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_501_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_501_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_501_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_501_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_501_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_502_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_502_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_502_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_502_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_502_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_502_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_502_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_502_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_502_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_502_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_502_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_502_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_502_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_502_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_502_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_503_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_503_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_503_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_503_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_503_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_503_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_503_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_503_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_503_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_503_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_503_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_503_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_503_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_503_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_503_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_503_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_503_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_504_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_504_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_504_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_504_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_504_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_504_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_504_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_504_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_504_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_504_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_504_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_504_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_504_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_504_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_504_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_504_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_504_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_504_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_504_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_504_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_504_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_504_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_504_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_504_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_504_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_504_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_504_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_504_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_505_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_505_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_505_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_505_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_505_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_505_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_505_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_505_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_505_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_505_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_505_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_505_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_505_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_506_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_506_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_506_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_506_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_506_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_506_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_506_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_506_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_506_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_506_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_506_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_506_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_506_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_506_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_506_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_506_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_506_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_506_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_506_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_506_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_506_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_506_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_506_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_507_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_507_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_507_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_507_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_507_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_507_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_507_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_507_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_507_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_507_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_507_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_507_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_507_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_507_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_507_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_507_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_507_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_508_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_508_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_508_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_508_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_508_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_508_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_508_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_508_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_508_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_508_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_509_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_509_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_509_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_509_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_509_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_509_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_509_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_509_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_509_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_509_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_509_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_510_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_510_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_510_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_511_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_511_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_511_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_511_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_511_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_511_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_511_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_511_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_511_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_512_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_512_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_512_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_512_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_512_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_512_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_512_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_512_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_512_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_512_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_512_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_513_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_513_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_513_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_513_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_513_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_513_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_513_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_513_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_513_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_513_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_514_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_514_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_514_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_514_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_514_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_514_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_514_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_515_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_515_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_515_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_515_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_515_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_515_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_515_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_515_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_515_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_515_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_515_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_515_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_515_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_516_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_516_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_516_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_516_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_516_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_516_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_516_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_516_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_516_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_516_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_516_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_516_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_516_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_516_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_517_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_517_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_517_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_517_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_517_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_517_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_517_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_517_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_517_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_517_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_517_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_517_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_517_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_517_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_517_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_518_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_518_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_518_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_518_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_518_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_518_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_518_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_518_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_518_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_518_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_519_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_519_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_519_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_519_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_519_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_519_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_519_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_519_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_519_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_519_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_519_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_520_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_520_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_520_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_520_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_520_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_520_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_520_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_520_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_520_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_520_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_520_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_520_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_520_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_520_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_521_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_521_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_521_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_521_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_521_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_521_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_522_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_522_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_522_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_522_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_522_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_522_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_522_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_522_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_522_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_522_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_522_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_522_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_522_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_522_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_523_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_523_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_523_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_523_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_523_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_523_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_524_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_524_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_524_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_524_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_524_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_524_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_524_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_524_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_524_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_524_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_524_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_524_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_524_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_524_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_524_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_524_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_524_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_524_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_524_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_524_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_524_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_524_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_524_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_524_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_524_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_525_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_525_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_525_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_525_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_525_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_525_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_525_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_525_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_525_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_525_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_525_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_525_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_525_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_525_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_525_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_525_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_525_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_525_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_525_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_525_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_525_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_525_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_525_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_526_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_526_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_526_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_526_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_526_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_526_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_526_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_526_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_526_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_526_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_526_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_526_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_526_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_526_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_526_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_526_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_526_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_526_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_526_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_527_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_527_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_527_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_527_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_527_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_527_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_527_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_527_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_527_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_527_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_527_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_527_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_527_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_527_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_527_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_527_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_527_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_527_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_528_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_528_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_528_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_528_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_528_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_528_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_528_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_528_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_528_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_528_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_528_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_528_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_529_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_529_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_529_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_529_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_529_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_529_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_529_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_529_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_529_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_529_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_529_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_529_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_529_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_529_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_529_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_529_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_529_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_529_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_529_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_529_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_529_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_529_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_530_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_530_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_530_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_530_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_530_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_530_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_530_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_530_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_530_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_530_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_530_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_530_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_530_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_530_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_531_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_531_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_531_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_531_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_531_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_531_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_531_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_531_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_531_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_531_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_531_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_531_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_532_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_532_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_532_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_532_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_532_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_532_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_532_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_532_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_532_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_532_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_532_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_532_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_532_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_532_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_532_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_532_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_532_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_532_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_532_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_532_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_532_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_532_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_532_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_532_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_532_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_533_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_533_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_533_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_533_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_533_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_533_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_533_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_533_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_533_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_534_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_534_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_534_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_534_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_534_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_534_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_534_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_534_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_534_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_534_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_534_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_534_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_534_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_534_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_534_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_534_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_534_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_535_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_535_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_535_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_535_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_535_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_535_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_535_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_535_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_535_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_535_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_535_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_535_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_535_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_535_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_535_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_535_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_535_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_535_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_535_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_536_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_536_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_536_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_536_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_536_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_536_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_536_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_536_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_536_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_536_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_536_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_536_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_536_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_536_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_536_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_536_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_536_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_536_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_536_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_536_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_536_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_536_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_536_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_536_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_536_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_536_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_537_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_537_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_537_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_537_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_537_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_537_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_537_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_537_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_537_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_537_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_537_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_537_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_537_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_537_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_537_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_537_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_537_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_537_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_538_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_538_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_538_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_538_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_538_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_538_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_538_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_538_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_538_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_538_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_538_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_538_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_538_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_538_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_538_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_538_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_538_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_538_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_539_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_539_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_539_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_539_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_539_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_539_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_539_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_540_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_540_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_540_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_540_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_540_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_540_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_540_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_540_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_540_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_540_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_540_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_540_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_540_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_541_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_541_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_541_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_541_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_541_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_541_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_541_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_541_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_542_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_542_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_542_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_542_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_542_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_542_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_542_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_542_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_542_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_542_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_542_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_542_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_542_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_542_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_542_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_542_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_542_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_542_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_542_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_542_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_542_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_542_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_542_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_542_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_543_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_543_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_543_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_543_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_543_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_543_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_543_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_543_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_543_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_543_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_543_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_543_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_543_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_543_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_543_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_543_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_544_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_544_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_544_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_544_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_544_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_544_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_544_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_544_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_544_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_544_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_544_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_544_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_544_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_544_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_544_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_544_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_544_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_544_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_544_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_545_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_545_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_545_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_545_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_545_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_545_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_545_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_546_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_546_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_546_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_546_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_546_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_546_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_546_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_546_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_546_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_546_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_546_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_546_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_546_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_546_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_546_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_547_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_547_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_547_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_547_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_547_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_547_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_547_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_547_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_547_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_547_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_547_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_547_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_547_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_547_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_547_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_547_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_547_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_548_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_548_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_548_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_548_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_548_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_548_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_548_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_548_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_548_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_548_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_548_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_548_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_548_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_548_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_548_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_548_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_548_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_549_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_549_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_549_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_549_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_549_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_549_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_549_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_549_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_549_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_550_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_550_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_550_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_550_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_550_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_550_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_550_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_550_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_550_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_550_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_550_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_550_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_550_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_550_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_550_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_550_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_550_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_551_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_551_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_551_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_551_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_551_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_551_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_552_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_552_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_552_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_552_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_552_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_552_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_552_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_552_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_552_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_552_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_552_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_552_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_552_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_552_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_552_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_552_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_553_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_553_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_553_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_553_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_553_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_553_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_553_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_553_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_553_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_553_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_553_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_553_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_553_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_553_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_553_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_553_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_553_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_554_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_554_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_554_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_554_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_554_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_554_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_554_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_554_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_554_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_554_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_554_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_554_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_554_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_554_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_554_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_554_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_554_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_554_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_554_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_555_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_555_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_555_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_555_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_555_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_555_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_555_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_555_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_555_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_555_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_555_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_555_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_556_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_556_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_556_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_556_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_556_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_556_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_556_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_556_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_556_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_556_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_556_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_556_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_556_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_556_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_556_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_556_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_557_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_557_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_557_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_557_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_557_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_557_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_557_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_557_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_557_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_557_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_557_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_557_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_557_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_557_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_557_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_557_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_557_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_557_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_557_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_557_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_558_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_558_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_558_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_558_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_558_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_558_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_558_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_558_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_558_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_558_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_558_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_558_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_558_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_558_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_558_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_558_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_558_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_558_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_558_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_558_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_558_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_558_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_558_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_559_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_559_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_559_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_559_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_559_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_559_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_559_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_559_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_559_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_559_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_559_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_559_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_560_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_560_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_560_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_560_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_560_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_560_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_560_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_560_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_560_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_560_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_560_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_560_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_560_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_560_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_560_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_560_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_560_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_560_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_560_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_560_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_560_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_561_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_561_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_561_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_561_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_561_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_561_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_562_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_562_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_562_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_562_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_562_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_562_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_562_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_562_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_562_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_562_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_562_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_562_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_562_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_562_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_562_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_562_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_562_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_562_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_562_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_562_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_562_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_562_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_562_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_562_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_562_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_563_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_563_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_563_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_563_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_563_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_563_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_563_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_563_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_563_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_563_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_563_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_563_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_563_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_563_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_563_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_563_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_563_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_563_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_563_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_563_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_563_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_563_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_563_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_563_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_563_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_563_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_563_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_563_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_564_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_564_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_564_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_564_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_564_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_564_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_564_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_564_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_564_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_564_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_564_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_564_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_564_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_564_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_564_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_564_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_564_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_564_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_564_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_564_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_564_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_564_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_564_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_565_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_565_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_565_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_565_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_565_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_565_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_565_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_565_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_565_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_566_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_566_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_566_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_566_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_566_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_566_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_566_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_566_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_566_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_566_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_566_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_566_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_566_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_566_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_566_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_566_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_566_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_567_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_567_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_567_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_567_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_567_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_567_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_567_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_567_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_567_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_567_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_567_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_567_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_567_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_567_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_567_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_568_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_568_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_568_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_568_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_568_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_568_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_568_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_568_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_568_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_568_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_568_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_568_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_568_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_568_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_568_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_568_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_568_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_568_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_568_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_568_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_568_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_568_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_568_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_569_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_569_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_569_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_569_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_569_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_569_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_569_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_569_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_569_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_569_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_569_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_570_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_570_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_570_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_570_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_570_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_570_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_570_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_570_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_570_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_570_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_570_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_570_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_570_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_570_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_570_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_570_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_571_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_571_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_571_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_571_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_571_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_571_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_571_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_571_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_572_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_572_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_572_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_572_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_572_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_572_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_572_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_572_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_572_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_572_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_572_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_572_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_572_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_572_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_572_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_572_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_572_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_572_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_572_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_573_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_573_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_573_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_573_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_573_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_573_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_573_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_573_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_573_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_573_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_573_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_574_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_574_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_574_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_574_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_574_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_574_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_574_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_574_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_574_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_574_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_574_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_574_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_574_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_574_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_574_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_574_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_574_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_574_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_574_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_575_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_575_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_575_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_575_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_575_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_575_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_575_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_575_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_575_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_575_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_575_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_575_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_575_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_575_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_575_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_575_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_575_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_575_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_575_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_575_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_576_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_576_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_576_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_576_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_576_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_576_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_576_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_576_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_576_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_576_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_576_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_576_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_576_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_576_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_576_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_576_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_577_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_577_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_577_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_577_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_577_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_577_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_577_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_577_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_577_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_578_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_578_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_578_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_578_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_578_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_578_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_578_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_578_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_578_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_578_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_578_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_578_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_578_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_579_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_579_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_579_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_579_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_579_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_579_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_579_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_579_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_579_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_579_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_579_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_579_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_579_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_579_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_579_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_579_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_579_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_579_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_580_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_580_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_580_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_580_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_580_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_580_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_580_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_580_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_580_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_580_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_580_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_580_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_580_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_580_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_580_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_580_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_580_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_580_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_580_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_580_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_580_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_580_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_580_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_580_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_580_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_581_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_581_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_581_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_581_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_581_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_581_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_581_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_581_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_581_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_581_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_581_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_581_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_581_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_581_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_581_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_582_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_582_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_582_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_582_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_582_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_582_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_582_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_582_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_582_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_582_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_582_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_582_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_582_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_582_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_582_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_582_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_582_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_583_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_583_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_583_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_583_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_583_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_583_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_583_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_583_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_583_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_583_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_583_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_583_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_583_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_583_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_583_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_583_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_583_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_584_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_584_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_584_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_584_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_584_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_584_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_584_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_584_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_584_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_584_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_585_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_585_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_585_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_585_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_585_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_585_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_585_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_585_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_586_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_586_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_586_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_586_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_586_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_586_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_586_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_586_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_586_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_586_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_586_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_586_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_586_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_586_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_586_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_586_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_586_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_587_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_587_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_587_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_587_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_587_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_587_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_587_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_587_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_587_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_587_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_587_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_587_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_587_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_587_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_588_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_588_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_588_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_588_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_588_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_588_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_588_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_588_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_588_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_588_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_588_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_588_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_588_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_588_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_588_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_588_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_589_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_589_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_589_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_590_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_590_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_590_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_590_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_590_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_590_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_590_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_590_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_590_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_590_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_590_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_590_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_590_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_590_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_591_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_591_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_591_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_591_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_591_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_591_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_591_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_591_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_591_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_591_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_591_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_591_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_591_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_591_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_591_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_592_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_592_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_592_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_592_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_592_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_592_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_592_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_592_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_592_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_592_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_592_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_592_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_592_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_592_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_592_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_592_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_592_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_592_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_592_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_592_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_592_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_592_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_593_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_593_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_593_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_593_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_593_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_593_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_593_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_593_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_593_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_593_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_593_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_593_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_593_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_593_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_593_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_593_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_593_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_593_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_593_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_593_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_593_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_593_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_593_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_593_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_593_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_593_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_594_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_594_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_594_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_594_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_594_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_594_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_594_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_594_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_594_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_594_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_594_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_594_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_594_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_594_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_594_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_594_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_594_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_594_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_594_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_594_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_594_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_594_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_595_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_595_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_595_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_595_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_595_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_595_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_595_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_595_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_595_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_595_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_595_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_595_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_595_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_595_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_595_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_595_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_595_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_596_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_596_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_596_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_596_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_596_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_596_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_596_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_596_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_596_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_596_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_596_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_596_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_596_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_596_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_596_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_596_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_596_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_596_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_596_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_596_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_597_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_597_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_597_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_597_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_597_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_597_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_597_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_597_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_597_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_597_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_597_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_597_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_597_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_597_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_597_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_597_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_597_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_598_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_598_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_598_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_598_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_598_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_598_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_598_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_598_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_598_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_598_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_598_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_598_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_599_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_599_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_599_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_599_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_599_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_599_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_599_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_599_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_599_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_599_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_599_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_599_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_599_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_600_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_600_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_600_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_600_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_600_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_600_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_600_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_600_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_600_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_600_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_600_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_600_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_600_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_600_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_600_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_601_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_601_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_601_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_601_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_601_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_601_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_601_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_601_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_602_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_602_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_602_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_602_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_602_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_602_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_602_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_602_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_602_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_602_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_602_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_602_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_602_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_603_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_603_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_603_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_603_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_603_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_603_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_603_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_603_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_603_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_603_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_603_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_603_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_603_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_603_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_603_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_603_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_603_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_603_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_603_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_604_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_604_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_604_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_604_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_604_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_604_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_604_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_604_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_604_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_604_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_604_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_604_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_604_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_604_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_604_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_604_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_604_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_604_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_604_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_605_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_605_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_605_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_605_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_605_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_605_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_605_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_605_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_605_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_605_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_605_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_605_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_605_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_605_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_605_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_605_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_605_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_605_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_605_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_605_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_606_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_606_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_606_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_606_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_606_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_606_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_606_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_606_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_606_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_606_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_606_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_606_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_606_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_606_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_606_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_606_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_606_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_607_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_607_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_607_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_607_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_607_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_607_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_607_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_607_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_607_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_607_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_607_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_607_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_607_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_607_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_607_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_607_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_608_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_608_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_608_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_608_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_608_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_608_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_608_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_608_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_608_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_608_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_608_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_608_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_608_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_608_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_608_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_608_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_608_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_608_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_608_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_608_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_608_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_609_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_609_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_609_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_609_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_609_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_609_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_609_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_609_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_609_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_609_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_609_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_609_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_609_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_609_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_609_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_609_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_609_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_609_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_609_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_610_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_610_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_610_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_610_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_610_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_610_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_610_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_610_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_610_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_610_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_610_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_610_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_610_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_611_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_611_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_611_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_611_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_611_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_611_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_611_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_611_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_611_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_611_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_611_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_611_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_611_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_611_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_611_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_611_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_612_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_612_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_612_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_612_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_612_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_612_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_612_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_612_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_612_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_612_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_612_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_612_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_612_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_612_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_612_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_612_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_612_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_612_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_612_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_613_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_613_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_613_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_613_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_613_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_613_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_613_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_613_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_613_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_613_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_613_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_613_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_613_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_613_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_613_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_613_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_614_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_614_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_614_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_614_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_614_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_614_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_614_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_614_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_614_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_614_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_614_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_614_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_614_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_615_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_615_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_615_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_615_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_615_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_615_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_615_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_615_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_615_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_615_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_615_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_616_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_616_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_616_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_616_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_616_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_616_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_616_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_616_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_616_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_616_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_616_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_616_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_616_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_616_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_616_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_616_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_616_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_616_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_617_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_617_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_617_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_617_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_617_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_617_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_617_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_618_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_618_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_618_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_618_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_618_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_618_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_618_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_618_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_618_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_618_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_618_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_618_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_618_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_618_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_618_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_618_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_619_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_619_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_619_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_619_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_619_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_619_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_619_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_619_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_619_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_619_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_619_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_619_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_619_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_619_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_619_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_619_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_619_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_619_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_619_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_619_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_619_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_620_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_620_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_620_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_620_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_620_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_620_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_620_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_620_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_620_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_620_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_620_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_620_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_620_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_620_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_620_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_620_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_620_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_620_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_620_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_620_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_620_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_621_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_621_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_621_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_621_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_621_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_621_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_621_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_621_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_622_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_622_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_622_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_622_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_622_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_622_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_622_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_622_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_622_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_622_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_622_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_622_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_622_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_622_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_622_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_622_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_622_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_622_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_623_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_623_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_623_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_623_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_623_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_623_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_623_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_623_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_623_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_623_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_623_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_623_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_623_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_623_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_623_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_624_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_624_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_624_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_624_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_624_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_624_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_624_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_624_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_624_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_624_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_624_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_624_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_624_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_624_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_624_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_624_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_624_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_624_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_624_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_625_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_625_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_625_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_625_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_625_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_625_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_625_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_625_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_625_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_625_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_626_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_626_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_626_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_626_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_626_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_626_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_626_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_626_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_626_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_626_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_626_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_626_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_626_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_626_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_626_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_626_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_627_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_627_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_627_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_627_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_627_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_627_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_627_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_627_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_627_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_627_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_627_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_627_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_627_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_627_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_627_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_627_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_627_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_627_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_627_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_627_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_627_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_627_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_628_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_628_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_628_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_628_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_628_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_628_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_628_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_628_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_628_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_628_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_629_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_629_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_629_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_629_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_629_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_629_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_629_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_629_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_629_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_630_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_630_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_630_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_630_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_630_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_630_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_630_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_630_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_630_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_630_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_630_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_630_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_630_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_630_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_630_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_631_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_631_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_631_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_631_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_631_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_631_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_631_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_631_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_631_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_631_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_631_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_631_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_631_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_631_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_631_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_631_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_632_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_632_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_632_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_632_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_632_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_632_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_632_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_632_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_632_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_632_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_632_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_632_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_632_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_632_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_632_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_632_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_632_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_632_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_632_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_632_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_632_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_632_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_632_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_632_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_632_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_633_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_633_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_633_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_633_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_633_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_633_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_633_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_633_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_633_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_633_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_634_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_634_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_634_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_634_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_634_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_634_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_634_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_634_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_634_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_634_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_634_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_634_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_634_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_634_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_634_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_634_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_634_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_634_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_634_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_634_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_635_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_635_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_635_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_635_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_635_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_635_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_635_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_635_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_635_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_635_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_635_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_635_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_635_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_635_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_635_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_635_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_635_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_636_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_636_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_636_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_636_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_636_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_636_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_636_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_636_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_636_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_636_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_636_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_636_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_636_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_636_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_636_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_636_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_637_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_637_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_637_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_637_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_637_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_637_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_637_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_637_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_637_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_637_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_637_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_637_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_637_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_637_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_637_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_637_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_637_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_637_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_638_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_638_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_638_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_638_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_638_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_638_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_638_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_638_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_638_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_638_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_638_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_638_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_638_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_638_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_638_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_638_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_638_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_638_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_639_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_639_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_639_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_639_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_639_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_639_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_639_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_639_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_639_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_640_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_640_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_640_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_640_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_640_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_640_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_640_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_640_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_640_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_640_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_640_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_640_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_640_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_640_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_640_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_640_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_640_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_640_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_640_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_641_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_641_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_641_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_641_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_641_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_641_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_641_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_641_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_641_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_641_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_641_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_641_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_641_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_641_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_642_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_642_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_642_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_642_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_642_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_642_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_642_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_642_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_642_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_642_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_642_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_642_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_642_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_642_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_642_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_642_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_642_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_643_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_643_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_643_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_643_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_643_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_643_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_643_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_643_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_643_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_643_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_643_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_644_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_644_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_644_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_644_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_644_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_644_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_644_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_644_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_644_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_644_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_644_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_644_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_644_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_644_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_644_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_644_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_644_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_644_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_644_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_644_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_645_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_645_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_645_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_645_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_645_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_645_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_645_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_645_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_645_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_645_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_645_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_645_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_645_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_645_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_645_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_646_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_646_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_646_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_646_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_646_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_646_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_646_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_646_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_646_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_646_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_646_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_646_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_646_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_646_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_646_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_646_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_646_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_646_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_646_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_646_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_646_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_646_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_646_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_646_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_646_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_647_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_647_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_647_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_647_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_647_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_647_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_647_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_647_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_647_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_647_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_647_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_647_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_647_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_647_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_647_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_647_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_647_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_647_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_647_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_648_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_648_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_648_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_648_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_648_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_648_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_648_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_648_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_648_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_648_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_648_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_648_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_648_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_648_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_648_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_648_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_648_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_648_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_648_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_648_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_648_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_648_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_648_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_648_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_648_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_648_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_649_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_649_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_649_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_649_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_649_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_649_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_649_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_649_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_649_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_649_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_649_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_649_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_649_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_649_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_649_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_649_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_649_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_649_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_649_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_649_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_650_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_650_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_650_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_650_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_650_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_650_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_650_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_650_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_650_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_650_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_650_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_650_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_650_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_650_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_651_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_651_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_651_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_651_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_651_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_651_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_651_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_651_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_651_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_651_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_652_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_652_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_652_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_652_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_652_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_652_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_652_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_652_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_652_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_652_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_652_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_652_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_652_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_653_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_653_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_653_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_653_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_653_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_653_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_653_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_653_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_653_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_653_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_653_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_653_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_653_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_653_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_654_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_654_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_654_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_654_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_654_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_654_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_654_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_654_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_654_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_654_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_654_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_654_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_654_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_654_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_654_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_654_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_654_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_654_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_654_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_655_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_655_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_655_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_655_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_655_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_655_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_655_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_655_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_655_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_655_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_655_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_655_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_655_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_656_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_656_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_656_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_656_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_656_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_656_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_656_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_656_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_656_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_656_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_656_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_656_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_656_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_656_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_656_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_656_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_656_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_656_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_656_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_656_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_656_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_656_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_656_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_656_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_657_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_657_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_657_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_657_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_657_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_657_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_657_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_657_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_657_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_657_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_657_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_657_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_657_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_657_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_657_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_657_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_657_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_658_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_658_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_658_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_658_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_658_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_658_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_658_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_658_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_658_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_658_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_658_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_658_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_658_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_658_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_659_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_659_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_659_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_659_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_659_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_659_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_659_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_659_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_659_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_659_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_659_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_660_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_660_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_660_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_660_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_660_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_660_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_660_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_660_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_660_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_660_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_661_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_661_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_661_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_661_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_661_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_661_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_661_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_661_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_661_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_661_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_661_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_661_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_661_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_661_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_662_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_662_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_662_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_662_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_662_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_662_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_662_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_662_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_662_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_662_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_662_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_662_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_662_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_662_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_662_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_662_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_662_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_662_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_663_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_663_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_663_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_663_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_663_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_663_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_663_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_663_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_663_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_663_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_663_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_663_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_663_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_663_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_663_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_663_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_663_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_663_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_663_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_663_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_663_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_664_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_664_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_664_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_664_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_664_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_664_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_664_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_664_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_664_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_664_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_664_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_664_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_664_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_664_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_664_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_664_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_664_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_664_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_664_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_665_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_665_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_665_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_665_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_665_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_665_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_665_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_665_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_665_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_665_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_665_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_665_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_665_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_665_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_666_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_666_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_666_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_666_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_667_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_667_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_667_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_667_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_667_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_667_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_667_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_667_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_667_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_667_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_667_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_667_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_667_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_667_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_668_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_668_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_668_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_668_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_668_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_668_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_668_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_668_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_668_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_668_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_668_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_668_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_668_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_668_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_668_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_668_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_669_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_669_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_669_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_669_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_669_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_669_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_669_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_669_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_669_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_669_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_669_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_670_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_670_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_670_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_670_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_670_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_670_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_670_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_670_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_671_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_671_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_671_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_671_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_671_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_671_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_671_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_671_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_671_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_671_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_671_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_671_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_671_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_672_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_672_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_672_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_672_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_672_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_672_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_672_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_672_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_672_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_672_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_672_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_672_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_672_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_672_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_673_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_673_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_673_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_673_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_673_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_673_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_673_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_673_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_674_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_674_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_674_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_674_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_674_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_674_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_674_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_674_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_675_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_675_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_675_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_675_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_675_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_675_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_675_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_675_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_675_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_675_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_675_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_675_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_675_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_675_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_675_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_675_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_676_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_676_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_676_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_676_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_676_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_676_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_676_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_676_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_676_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_676_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_676_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_676_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_676_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_676_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_676_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_677_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_677_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_677_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_677_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_677_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_677_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_677_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_677_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_677_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_677_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_678_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_678_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_678_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_678_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_678_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_678_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_678_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_678_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_678_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_678_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_678_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_678_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_678_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_678_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_678_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_679_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_679_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_680_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_680_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_680_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_680_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_680_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_680_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_680_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_680_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_681_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_681_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_681_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_681_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_681_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_681_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_681_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_681_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_681_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_681_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_681_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_681_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_681_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_681_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_681_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_681_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_682_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_682_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_682_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_682_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_682_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_682_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_682_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_682_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_682_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_683_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_683_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_683_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_683_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_683_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_683_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_683_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_683_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_683_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_683_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_683_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_683_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_683_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_683_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_683_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_683_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_684_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_684_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_684_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_684_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_684_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_684_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_684_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_684_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_685_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_685_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_686_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_686_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_687_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_687_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_687_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_687_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_687_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_687_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_687_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_687_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_687_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_687_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_687_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_687_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_687_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_687_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_687_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_687_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_688_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_688_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_688_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_688_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_688_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_688_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_688_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_688_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_688_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_688_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_688_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_688_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_688_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_688_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_688_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_689_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_689_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_689_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_689_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_689_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_689_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_689_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_689_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_689_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_690_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_690_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_690_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_690_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_690_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_690_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_690_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_690_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_690_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_690_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_690_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_690_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_690_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_690_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_690_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_691_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_691_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_691_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_691_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_691_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_691_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_691_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_691_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_691_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_691_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_692_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_692_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_692_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_692_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_692_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_692_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_692_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_692_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_692_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_692_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_692_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_692_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_692_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_692_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_692_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_693_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_693_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_693_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_694_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_694_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_694_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_694_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_694_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_694_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_694_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_694_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_695_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_695_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_695_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_695_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_695_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_695_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_695_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_695_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_695_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_696_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_696_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_696_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_696_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_696_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_696_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_696_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_696_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_696_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_696_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_696_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_696_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_696_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_696_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_696_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_697_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_697_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_697_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_697_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_697_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_697_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_697_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_697_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_697_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_697_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_697_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_697_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_697_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_697_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_697_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_697_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_698_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_698_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_698_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_698_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_698_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_698_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_698_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_698_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_698_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_698_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_698_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_698_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_698_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_698_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_698_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_699_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_699_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_699_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_699_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_699_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_699_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_699_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_699_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_699_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_700_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_700_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_700_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_700_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_700_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_700_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_700_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_700_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_700_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_700_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_700_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_700_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_700_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_700_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_700_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_701_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_701_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_702_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_702_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_702_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_702_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_702_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_702_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_702_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_702_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_702_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_702_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_702_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_702_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_702_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_702_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_702_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_703_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_703_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_703_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_703_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_703_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_703_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_703_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_703_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_703_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_703_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_703_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_703_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_703_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_703_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_703_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_703_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_704_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_704_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_704_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_704_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_704_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_704_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_704_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_704_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_704_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_704_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_704_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_704_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_704_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_704_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_704_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_705_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_705_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_705_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_705_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_705_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_705_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_705_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_705_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_705_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_707_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_707_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_707_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_707_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_707_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_707_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_707_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_707_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_708_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_708_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_708_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_708_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_708_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_708_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_708_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_708_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_708_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_708_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_708_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_708_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_708_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_708_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_708_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_709_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_709_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_709_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_709_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_709_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_709_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_709_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_709_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_710_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_710_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_710_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_710_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_710_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_710_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_710_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_710_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_710_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_710_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_710_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_710_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_710_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_710_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_710_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_711_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_711_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_711_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_711_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_711_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_711_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_711_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_711_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_712_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_712_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_712_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_712_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_712_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_712_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_712_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_712_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_713_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_713_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_713_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_713_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_713_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_713_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_713_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_713_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_713_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_713_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_713_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_713_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_713_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_713_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_713_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_714_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_714_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_714_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_714_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_714_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_714_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_714_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_714_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_714_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_715_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_715_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_715_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_715_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_715_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_715_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_715_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_715_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_715_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_715_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_715_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_716_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_716_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_716_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_716_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_716_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_716_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_716_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_716_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_716_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_716_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_716_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_716_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_716_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_716_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_716_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_717_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_717_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_717_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_717_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_717_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_717_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_717_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_717_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_717_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_717_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_717_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_717_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_717_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_717_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_717_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_717_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_718_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_718_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_718_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_718_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_718_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_718_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_718_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_718_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_718_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_718_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_718_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_718_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_718_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_718_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_718_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_719_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_719_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_719_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_719_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_719_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_719_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_719_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_719_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_719_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_720_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_720_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_720_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_720_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_720_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_720_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_720_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_720_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_720_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_720_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_720_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_720_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_720_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_720_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_720_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_721_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_721_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_721_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_721_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_721_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_721_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_721_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_721_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_721_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_721_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_722_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_722_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_722_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_722_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_722_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_722_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_722_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_722_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_722_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_723_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_723_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_723_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_723_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_723_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_723_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_723_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_723_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_723_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_723_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_723_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_723_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_723_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_723_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_723_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_724_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_724_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_724_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_724_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_724_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_724_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_724_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_724_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_724_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_724_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_724_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_724_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_724_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_724_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_724_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_725_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_725_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_725_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_725_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_725_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_725_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_725_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_725_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_725_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_726_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_726_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_726_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_726_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_726_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_726_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_726_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_726_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_726_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_726_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_726_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_726_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_726_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_726_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_726_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_727_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_727_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_727_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_727_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_727_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_727_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_727_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_727_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_727_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_728_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_728_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_728_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_728_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_728_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_728_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_728_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_728_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_729_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_729_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_729_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_729_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_729_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_729_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_729_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_730_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_730_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_730_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_730_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_730_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_730_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_730_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_730_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_730_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_730_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_730_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_730_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_730_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_730_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_730_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_731_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_731_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_731_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_731_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_731_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_731_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_731_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_731_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_731_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_731_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_731_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_731_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_731_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_731_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_731_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_731_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_732_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_732_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_732_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_732_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_732_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_732_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_732_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_732_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_732_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_732_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_732_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_732_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_732_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_732_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_732_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_733_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_733_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_733_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_733_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_733_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_733_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_733_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_733_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_733_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_733_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_733_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_733_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_733_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_733_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_733_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_733_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_734_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_734_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_734_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_734_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_734_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_734_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_734_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_734_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_734_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_734_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_734_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_734_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_734_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_734_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_735_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_735_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_735_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_735_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_735_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_735_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_735_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_735_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_735_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_736_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_736_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_736_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_736_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_736_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_736_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_736_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_736_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_736_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_736_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_736_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_736_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_736_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_736_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_736_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_737_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_737_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_737_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_737_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_737_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_737_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_737_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_737_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_738_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_738_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_738_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_738_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_738_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_738_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_738_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_738_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_739_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_739_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_739_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_739_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_739_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_739_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_739_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_739_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_739_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_739_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_739_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_739_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_739_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_739_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_739_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_740_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_740_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_740_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_741_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_741_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_741_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_741_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_741_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_741_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_741_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_741_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_742_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_742_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_742_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_742_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_742_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_742_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_742_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_742_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_742_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_742_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_742_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_742_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_742_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_742_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_742_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_743_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_743_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_743_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_743_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_743_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_743_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_743_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_743_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_743_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_743_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_743_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_743_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_743_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_743_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_743_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_743_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_744_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_744_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_744_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_744_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_744_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_744_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_744_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_744_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_744_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_744_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_744_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_744_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_744_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_744_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_744_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_745_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_745_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_745_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_745_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_745_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_745_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_745_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_745_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_745_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_745_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_746_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_746_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_746_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_746_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_746_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_746_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_746_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_746_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_746_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_747_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_747_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_747_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_747_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_747_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_747_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_747_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_747_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_747_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_747_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_747_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_747_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_747_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_747_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_747_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_747_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_748_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_748_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_748_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_748_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_748_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_748_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_748_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_748_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_748_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_748_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_748_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_748_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_748_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_748_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_748_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_749_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_749_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_749_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_750_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_750_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_750_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_750_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_750_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_750_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_750_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_750_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_751_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_751_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_751_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_751_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_751_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_751_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_751_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_751_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_751_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_752_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_752_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_752_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_752_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_752_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_752_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_752_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_752_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_752_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_752_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_752_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_752_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_752_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_752_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_752_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_753_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_753_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_753_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_753_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_753_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_753_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_753_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_753_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_753_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_753_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_753_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_753_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_753_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_753_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_753_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_753_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_754_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_754_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_754_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_754_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_754_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_754_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_754_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_754_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_755_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_755_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_755_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_755_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_755_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_755_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_755_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_755_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_755_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_756_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_756_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_756_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_756_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_756_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_756_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_756_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_756_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_756_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_756_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_756_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_756_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_756_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_756_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_756_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_757_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_758_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_758_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_758_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_758_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_758_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_758_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_758_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_758_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_758_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_758_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_758_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_758_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_758_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_758_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_758_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_759_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_759_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_759_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_759_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_759_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_759_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_759_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_759_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_759_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_759_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_759_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_759_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_759_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_759_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_759_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_759_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_760_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_760_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_760_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_760_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_760_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_760_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_760_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_760_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_760_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_760_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_760_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_760_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_760_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_760_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_760_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_761_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_761_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_761_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_761_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_761_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_761_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_761_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_761_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_761_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_762_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_762_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_762_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_762_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_762_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_762_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_762_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_762_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_762_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_762_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_762_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_762_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_762_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_762_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_762_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_763_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_763_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_763_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_763_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_763_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_763_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_763_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_763_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_763_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_764_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_764_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_764_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_764_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_764_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_764_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_764_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_764_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_764_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_764_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_764_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_764_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_764_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_764_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_765_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_765_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_765_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_765_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_765_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_765_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_765_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_765_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_765_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_765_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_765_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_765_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_765_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_765_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_765_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_765_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_766_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_766_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_766_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_766_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_766_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_766_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_766_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_766_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_766_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_766_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_766_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_766_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_766_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_766_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_766_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_767_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_767_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_767_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_767_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_767_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_767_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_767_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_767_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_767_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_767_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_767_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_767_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_767_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_767_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_767_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_768_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_768_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_768_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_768_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_768_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_768_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_768_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_768_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_768_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_768_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_768_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_768_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_768_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_768_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_769_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_769_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_769_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_769_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_769_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_769_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_769_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_769_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_769_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_770_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_770_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_770_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_770_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_770_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_770_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_770_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_771_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_771_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_771_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_771_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_771_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_771_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_771_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_771_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_771_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_771_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_772_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_772_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_772_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_772_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_772_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_772_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_772_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_772_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_772_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_772_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_772_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_772_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_772_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_772_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_772_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_773_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_773_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_773_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_773_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_773_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_773_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_773_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_773_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_773_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_773_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_774_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_774_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_774_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_774_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_774_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_774_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_774_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_774_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_774_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_775_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_775_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_775_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_775_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_775_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_775_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_775_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_775_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_775_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_775_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_775_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_775_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_775_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_775_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_775_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_775_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_776_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_776_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_776_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_776_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_776_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_776_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_776_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_776_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_776_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_776_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_776_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_776_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_776_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_776_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_776_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_777_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_777_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_777_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_777_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_777_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_777_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_777_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_777_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_777_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_777_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_777_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_777_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_777_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_777_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_777_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_777_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_778_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_778_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_778_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_778_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_778_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_778_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_778_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_778_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_778_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_779_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_779_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_779_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_779_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_779_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_779_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_779_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_779_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_780_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_780_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_780_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_780_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_780_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_780_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_780_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_780_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_780_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_780_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_780_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_780_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_780_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_780_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_780_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_781_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_781_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_781_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_781_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_781_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_781_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_781_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_781_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_781_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_781_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_781_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_781_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_781_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_781_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_781_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_781_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_782_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_782_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_782_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_782_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_782_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_782_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_782_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_782_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_782_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_782_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_782_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_782_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_782_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_782_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_782_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_783_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_783_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_783_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_783_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_783_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_783_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_783_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_783_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_783_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_784_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_784_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_784_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_784_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_784_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_784_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_784_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_784_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_784_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_784_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_784_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_784_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_784_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_784_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_784_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_785_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_785_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_785_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_785_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_785_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_785_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_785_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_785_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_786_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_786_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_786_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_786_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_786_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_786_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_786_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_786_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_786_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_786_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_786_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_786_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_786_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_786_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_786_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_787_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_787_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_787_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_787_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_787_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_787_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_787_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_787_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_787_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_787_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_787_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_787_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_787_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_787_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_787_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_788_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_788_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_788_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_788_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_788_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_788_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_788_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_788_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_788_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_788_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_788_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_788_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_788_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_788_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_788_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_789_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_789_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_789_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_789_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_789_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_789_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_789_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_789_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_789_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_789_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_789_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_789_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_789_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_789_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_789_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_789_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_790_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_790_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_790_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_790_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_790_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_790_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_790_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_790_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_790_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_790_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_790_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_790_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_790_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_790_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_790_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_791_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_791_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_791_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_791_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_791_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_791_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_791_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_791_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_791_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_791_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_791_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_791_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_791_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_791_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_791_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_792_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_792_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_792_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_792_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_792_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_792_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_792_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_792_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_793_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_793_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_793_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_793_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_793_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_793_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_793_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_793_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_793_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_793_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_793_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_793_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_793_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_793_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_793_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_793_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_794_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_794_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_794_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_794_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_794_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_794_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_794_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_794_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_795_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_795_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_795_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_795_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_795_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_795_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_795_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_795_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_795_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_796_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_796_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_796_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_796_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_796_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_796_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_796_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_796_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_796_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_796_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_796_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_796_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_796_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_796_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_796_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_797_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_797_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_797_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_797_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_797_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_797_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_797_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_797_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_797_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_797_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_797_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_797_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_797_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_797_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_797_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_798_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_798_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_798_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_798_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_798_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_798_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_798_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_798_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_799_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_799_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_799_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_799_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_799_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_799_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_799_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_799_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_799_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_799_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_800_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_800_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_800_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_800_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_800_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_800_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_800_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_800_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_800_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_800_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_800_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_800_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_800_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_800_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_800_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_801_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_801_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_801_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_801_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_801_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_801_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_801_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_801_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_801_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_801_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_801_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_801_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_801_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_801_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_801_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_801_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_802_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_802_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_802_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_802_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_802_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_802_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_802_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_802_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_802_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_803_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_803_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_803_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_803_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_803_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_803_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_803_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_803_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_803_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_803_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_803_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_803_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_803_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_803_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_803_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_803_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_804_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_804_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_804_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_804_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_804_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_804_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_804_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_804_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_804_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_804_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_804_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_804_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_804_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_804_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_804_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_805_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_805_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_805_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_805_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_805_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_805_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_805_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_805_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_805_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_806_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_806_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_806_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_806_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_806_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_806_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_806_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_806_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_807_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_807_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_807_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_807_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_807_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_807_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_807_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_807_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_807_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_808_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_808_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_808_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_808_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_808_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_808_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_808_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_808_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_808_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_808_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_808_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_808_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_808_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_808_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_808_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_809_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_809_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_809_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_809_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_809_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_809_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_809_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_809_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_809_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_810_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_810_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_810_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_810_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_810_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_810_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_810_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_810_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_810_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_810_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_810_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_810_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_810_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_810_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_810_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_811_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_811_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_811_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_811_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_811_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_811_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_811_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_811_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_811_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_812_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_812_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_812_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_812_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_812_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_812_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_812_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_812_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_812_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_812_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_812_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_812_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_812_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_812_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_812_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_813_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_813_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_813_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_813_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_813_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_813_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_813_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_813_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_814_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_814_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_814_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_814_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_814_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_814_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_814_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_814_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_814_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_815_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_815_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_815_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_815_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_815_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_815_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_815_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_815_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_815_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_815_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_816_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_816_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_816_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_816_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_816_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_816_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_816_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_816_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_816_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_816_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_816_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_816_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_816_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_816_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_816_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_817_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_817_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_817_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_817_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_817_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_817_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_817_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_817_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_817_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_818_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_818_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_818_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_818_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_818_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_818_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_818_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_818_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_819_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_819_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_819_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_819_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_819_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_819_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_819_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_819_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_819_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_819_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_820_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_820_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_820_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_820_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_820_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_820_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_820_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_820_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_820_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_820_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_820_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_820_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_820_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_820_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_820_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_821_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_821_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_821_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_821_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_821_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_821_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_821_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_821_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_821_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_821_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_822_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_822_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_822_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_822_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_822_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_822_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_822_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_822_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_822_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_822_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_822_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_822_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_822_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_822_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_823_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_823_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_823_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_823_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_823_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_823_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_823_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_823_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_823_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_823_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_823_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_823_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_823_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_823_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_823_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_824_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_824_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_824_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_824_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_824_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_824_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_824_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_824_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_824_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_824_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_824_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_824_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_824_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_824_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_824_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_825_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_825_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_825_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_825_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_825_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_825_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_825_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_825_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_826_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_826_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_826_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_826_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_826_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_826_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_826_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_826_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_826_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_826_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_826_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_826_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_826_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_826_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_826_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_827_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_827_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_827_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_827_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_827_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_827_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_827_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_827_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_827_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_827_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_827_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_827_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_827_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_827_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_827_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_827_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_828_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_828_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_828_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_828_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_828_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_828_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_828_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_828_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_828_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_829_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_829_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_829_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_829_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_829_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_829_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_829_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_829_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_829_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_829_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_829_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_829_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_829_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_829_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_829_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_829_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_830_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_830_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_830_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_830_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_830_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_830_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_830_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_830_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_830_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_830_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_830_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_830_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_830_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_830_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_830_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_831_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_831_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_831_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_831_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_831_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_831_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_831_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_831_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_831_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_831_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_831_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_831_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_831_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_831_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_831_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_831_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_832_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_832_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_832_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_832_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_832_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_832_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_832_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_832_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_832_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_832_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_832_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_832_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_832_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_832_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_832_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_833_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_833_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_833_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_833_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_833_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_833_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_833_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_833_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_833_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_833_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_833_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_833_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_833_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_833_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_833_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_833_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_834_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_834_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_835_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_835_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_835_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_835_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_835_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_835_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_835_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_835_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_835_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_835_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_835_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_835_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_835_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_835_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_835_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_836_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_836_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_836_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_836_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_836_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_836_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_836_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_836_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_836_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_837_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_837_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_837_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_837_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_837_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_837_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_837_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_837_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_837_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_837_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_837_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_837_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_837_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_837_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_837_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_837_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_838_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_838_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_838_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_838_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_838_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_838_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_838_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_838_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_838_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_838_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_838_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_838_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_838_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_838_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_838_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_839_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_839_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_839_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_839_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_839_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_839_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_839_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_839_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_839_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_840_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_840_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_840_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_840_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_840_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_840_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_840_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_840_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_840_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_840_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_840_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_840_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_840_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_840_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_840_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_841_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_841_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_841_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_841_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_841_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_841_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_841_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_842_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_842_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_842_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_842_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_842_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_842_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_842_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_842_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_842_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_842_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_842_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_842_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_842_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_842_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_842_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_843_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_843_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_843_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_843_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_843_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_843_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_843_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_843_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_843_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_843_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_843_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_843_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_843_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_843_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_843_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_843_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_844_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_844_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_844_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_844_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_844_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_844_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_844_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_844_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_844_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_844_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_844_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_844_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_844_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_844_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_844_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_845_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_845_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_845_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_845_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_845_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_845_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_845_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_845_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_845_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_846_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_846_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_846_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_846_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_846_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_846_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_846_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_847_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_847_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_847_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_847_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_847_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_847_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_847_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_847_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_847_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_847_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_847_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_847_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_847_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_847_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_847_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_847_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_848_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_848_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_848_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_848_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_848_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_848_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_848_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_848_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_848_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_849_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_849_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_849_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_849_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_849_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_849_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_849_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_849_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_850_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_850_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_850_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_850_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_850_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_850_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_850_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_850_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_850_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_850_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_850_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_850_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_850_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_850_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_850_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_851_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_851_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_851_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_851_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_851_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_851_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_851_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_851_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_851_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_851_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_851_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_851_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_851_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_851_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_851_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_852_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_852_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_852_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_852_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_852_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_852_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_852_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_852_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_852_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_853_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_853_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_853_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_853_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_853_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_853_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_853_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_853_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_853_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_853_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_853_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_853_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_853_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_853_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_853_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_854_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_854_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_854_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_854_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_854_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_854_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_854_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_854_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_854_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_854_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_854_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_854_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_854_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_854_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_854_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_855_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_855_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_855_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_855_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_855_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_855_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_855_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_855_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_855_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_855_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_856_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_856_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_856_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_856_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_856_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_856_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_856_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_856_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_856_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_856_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_856_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_856_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_856_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_856_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_857_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_857_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_857_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_857_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_857_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_857_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_857_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_857_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_857_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_857_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_857_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_857_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_857_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_857_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_857_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_857_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_858_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_858_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_858_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_858_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_858_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_858_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_858_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_858_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_858_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_858_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_858_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_858_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_858_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_858_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_858_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_859_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_859_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_859_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_859_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_859_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_859_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_859_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_859_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_859_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_859_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_859_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_859_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_859_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_859_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_859_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_859_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_860_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_860_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_860_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_860_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_860_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_860_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_860_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_860_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_860_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_860_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_860_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_860_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_860_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_860_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_860_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_861_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_861_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_861_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_861_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_861_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_861_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_861_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_861_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_861_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_861_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_862_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_862_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_862_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_862_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_862_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_862_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_862_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_862_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_862_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_862_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_862_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_862_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_862_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_862_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_862_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_863_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_863_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_863_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_863_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_863_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_863_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_863_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_863_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_863_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_863_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_864_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_864_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_864_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_864_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_864_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_864_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_864_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_864_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_864_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_864_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_864_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_864_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_864_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_864_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_864_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_865_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_865_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_865_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_865_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_865_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_865_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_865_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_865_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_865_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_865_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_865_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_865_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_865_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_865_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_865_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_865_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_866_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_866_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_866_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_866_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_866_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_866_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_866_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_866_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_866_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_866_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_866_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_866_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_866_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_866_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_866_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_867_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_867_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_867_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_867_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_867_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_867_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_867_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_867_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_867_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_868_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_868_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_868_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_868_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_868_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_868_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_868_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_868_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_868_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_868_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_868_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_868_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_868_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_868_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_868_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_869_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_869_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_869_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_869_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_869_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_869_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_869_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_870_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_870_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_870_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_870_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_870_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_870_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_870_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_870_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_870_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_870_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_870_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_870_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_870_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_870_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_870_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_871_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_871_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_871_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_871_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_871_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_871_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_871_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_871_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_871_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_871_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_871_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_871_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_871_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_871_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_871_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_871_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_872_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_872_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_872_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_872_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_872_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_872_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_872_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_872_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_872_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_873_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_873_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_873_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_874_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_874_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_874_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_874_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_874_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_874_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_874_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_874_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_874_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_874_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_874_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_874_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_874_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_874_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_874_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_875_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_875_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_875_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_875_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_875_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_875_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_875_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_875_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_875_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_875_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_875_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_876_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_876_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_876_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_876_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_876_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_876_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_876_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_876_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_876_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_876_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_876_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_876_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_876_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_876_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_877_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_877_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_877_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_877_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_877_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_877_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_877_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_877_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_877_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_877_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_877_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_877_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_877_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_877_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_877_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_877_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_878_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_878_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_878_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_878_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_878_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_878_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_878_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_878_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_878_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_878_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_878_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_878_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_878_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_878_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_878_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_879_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_879_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_879_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_879_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_879_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_879_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_879_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_879_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_880_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_880_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_880_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_880_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_880_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_880_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_880_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_880_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_880_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_880_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_880_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_880_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_880_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_880_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_881_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_881_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_881_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_881_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_881_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_881_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_881_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_881_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_882_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_882_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_882_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_882_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_882_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_882_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_882_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_882_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_882_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_883_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_883_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_883_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_883_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_883_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_883_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_883_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_883_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_883_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_883_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_883_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_883_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_883_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_883_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_883_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_883_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_884_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_884_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_884_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_884_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_884_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_884_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_884_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_884_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_884_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_885_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_885_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_885_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_885_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_885_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_885_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_885_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_885_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_885_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_885_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_885_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_885_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_885_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_885_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_885_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_885_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_886_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_886_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_886_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_886_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_886_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_886_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_886_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_886_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_886_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_887_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_887_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_887_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_887_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_887_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_887_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_887_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_887_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_887_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_887_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_887_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_887_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_887_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_887_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_887_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_887_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_888_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_888_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_888_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_888_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_888_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_888_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_888_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_888_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_888_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_888_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_888_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_888_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_888_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_888_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_888_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_889_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_889_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_889_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_889_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_889_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_889_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_889_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_889_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_889_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_889_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_890_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_890_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_890_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_890_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_890_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_890_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_890_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_890_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_890_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_890_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_890_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_890_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_890_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_890_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_890_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_891_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_891_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_891_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_891_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_891_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_891_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_891_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_891_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_891_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_892_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_892_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_892_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_892_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_892_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_892_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_892_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_892_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_892_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_892_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_892_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_892_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_892_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_892_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_892_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_893_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_893_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_893_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_893_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_893_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_893_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_893_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_893_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_893_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_894_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_894_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_894_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_894_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_894_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_894_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_894_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_894_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_894_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_894_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_894_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_894_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_894_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_894_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_894_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_895_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_895_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_895_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_895_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_895_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_895_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_895_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_895_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_895_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_896_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_896_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_896_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_896_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_896_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_896_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_896_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_896_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_896_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_897_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_898_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_898_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_898_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_898_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_898_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_898_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_898_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_898_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_898_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_898_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_898_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_898_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_898_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_898_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_898_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_899_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_899_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_899_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_899_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_899_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_899_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_899_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_899_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_899_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_900_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_900_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_900_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_900_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_900_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_900_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_900_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_900_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_900_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_900_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_900_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_900_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_900_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_900_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_900_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_901_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_901_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_901_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_901_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_901_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_901_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_901_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_901_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_901_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_902_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_902_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_902_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_902_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_902_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_902_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_902_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_902_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_902_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_903_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_903_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_903_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_903_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_903_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_903_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_903_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_903_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_903_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_903_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_903_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_903_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_903_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_903_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_903_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_903_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_904_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_904_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_904_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_904_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_904_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_904_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_904_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_904_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_905_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_905_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_905_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_905_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_905_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_905_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_905_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_905_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_905_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_905_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_905_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_905_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_905_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_905_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_905_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_906_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_906_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_906_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_906_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_906_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_906_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_906_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_906_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_906_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_906_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_906_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_906_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_906_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_906_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_907_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_907_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_907_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_907_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_907_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_907_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_907_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_907_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_907_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_907_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_907_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_907_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_907_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_907_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_907_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_908_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_908_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_908_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_908_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_908_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_908_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_908_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_908_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_908_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_908_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_908_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_908_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_908_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_908_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_909_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_909_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_909_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_909_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_909_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_909_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_909_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_909_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_909_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_910_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_910_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_910_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_910_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_910_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_910_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_910_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_910_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_910_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_911_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_911_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_911_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_911_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_911_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_911_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_911_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_911_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_911_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_912_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_912_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_912_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_912_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_912_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_912_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_912_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_912_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_912_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_912_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_912_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_912_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_912_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_912_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_912_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_913_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_913_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_913_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_913_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_913_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_913_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_913_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_913_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_913_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_913_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_913_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_913_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_913_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_913_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_913_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_913_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_914_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_914_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_914_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_914_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_914_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_914_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_914_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_914_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_914_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_914_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_914_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_914_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_914_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_914_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_914_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_915_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_915_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_915_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_915_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_915_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_915_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_915_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_915_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_915_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_916_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_916_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_916_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_916_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_916_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_916_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_916_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_916_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_916_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_916_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_916_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_916_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_916_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_916_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_916_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_917_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_917_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_917_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_917_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_917_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_917_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_917_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_917_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_917_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_917_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_918_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_918_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_918_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_918_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_918_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_918_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_918_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_918_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_919_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_919_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_919_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_919_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_919_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_919_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_919_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_919_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_919_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_919_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_919_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_919_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_919_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_919_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_919_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_919_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_920_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_920_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_920_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_920_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_920_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_920_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_920_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_920_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_920_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_920_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_920_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_920_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_920_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_920_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_920_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_921_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_921_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_921_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_921_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_921_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_921_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_921_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_921_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_921_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_921_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_921_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_921_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_921_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_921_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_921_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_921_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_922_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_922_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_922_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_922_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_922_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_922_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_922_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_922_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_923_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_923_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_923_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_923_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_923_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_923_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_923_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_923_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_923_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_924_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_924_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_924_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_924_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_924_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_924_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_924_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_924_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_924_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_924_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_924_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_924_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_924_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_924_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_924_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_925_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_925_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_925_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_925_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_925_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_925_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_925_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_925_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_926_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_926_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_926_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_926_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_926_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_926_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_926_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_926_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_927_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_927_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_927_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_927_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_927_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_927_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_927_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_927_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_927_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_927_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_927_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_927_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_927_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_927_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_927_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_927_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_928_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_928_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_928_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_928_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_928_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_928_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_928_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_928_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_928_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_928_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_928_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_928_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_928_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_928_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_928_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_929_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_929_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_929_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_929_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_929_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_929_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_929_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_929_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_930_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_930_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_930_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_930_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_930_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_930_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_930_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_930_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_930_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_930_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_930_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_930_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_930_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_930_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_930_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_931_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_931_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_931_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_931_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_931_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_931_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_931_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_931_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_931_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_931_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_931_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_931_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_931_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_931_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_931_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_931_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_932_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_932_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_932_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_932_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_932_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_932_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_932_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_932_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_932_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_933_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_933_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_933_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_933_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_933_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_933_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_933_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_933_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_933_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_933_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_933_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_933_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_933_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_933_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_933_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_933_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_934_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_934_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_934_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_934_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_934_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_934_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_934_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_934_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_934_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_935_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_935_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_935_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_935_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_935_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_935_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_935_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_935_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_935_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_935_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_935_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_935_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_935_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_935_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_935_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_935_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_936_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_936_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_936_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_936_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_936_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_936_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_936_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_936_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_936_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_937_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_937_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_937_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_937_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_937_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_937_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_937_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_937_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_938_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_938_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_938_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_938_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_938_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_938_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_938_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_938_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_938_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_939_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_939_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_939_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_939_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_939_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_939_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_939_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_939_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_939_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_940_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_940_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_940_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_940_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_940_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_940_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_940_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_940_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_940_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_940_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_940_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_940_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_940_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_940_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_941_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_941_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_941_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_941_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_941_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_941_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_941_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_941_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_941_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_941_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_941_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_941_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_941_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_941_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_941_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_941_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_942_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_942_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_942_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_942_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_942_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_942_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_942_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_942_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_942_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_942_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_942_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_942_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_942_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_942_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_942_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_943_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_943_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_943_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_943_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_943_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_943_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_943_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_943_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_943_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_943_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_943_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_943_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_943_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_943_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_943_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_943_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_944_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_944_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_944_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_944_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_944_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_944_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_944_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_944_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_944_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_944_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_944_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_944_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_944_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_944_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_944_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_945_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_945_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_945_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_945_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_945_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_945_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_945_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_945_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_945_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_945_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_946_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_946_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_946_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_946_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_946_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_946_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_946_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_946_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_946_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_946_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_946_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_946_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_946_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_946_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_946_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_947_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_947_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_947_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_947_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_947_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_947_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_947_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_947_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_947_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_947_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_947_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_947_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_947_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_947_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_947_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_947_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_948_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_948_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_948_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_948_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_948_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_948_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_948_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_948_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_948_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_948_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_948_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_948_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_948_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_948_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_948_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_949_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_949_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_949_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_949_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_949_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_949_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_949_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_949_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_949_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_949_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_949_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_949_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_949_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_949_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_949_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_949_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_950_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_950_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_950_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_950_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_950_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_950_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_950_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_950_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_950_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_950_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_950_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_950_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_950_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_950_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_950_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_951_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_951_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_951_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_951_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_951_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_951_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_951_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_951_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_951_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_952_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_952_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_952_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_952_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_952_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_952_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_952_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_952_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_952_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_952_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_952_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_952_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_952_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_952_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_952_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_953_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_953_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_953_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_953_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_953_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_953_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_953_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_953_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_954_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_954_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_954_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_954_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_954_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_954_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_954_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_954_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_954_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_954_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_954_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_954_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_954_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_954_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_954_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_955_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_955_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_955_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_955_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_955_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_955_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_955_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_955_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_955_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_955_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_955_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_955_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_955_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_955_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_955_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_955_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_956_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_956_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_956_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_956_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_956_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_956_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_956_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_956_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_956_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_957_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_957_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_957_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_957_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_957_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_957_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_957_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_957_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_957_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_957_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_957_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_957_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_957_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_957_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_957_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_957_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_958_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_958_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_958_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_958_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_958_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_958_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_958_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_958_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_958_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_958_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_958_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_958_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_958_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_958_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_959_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_959_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_959_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_959_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_959_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_959_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_959_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_959_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_959_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_959_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_960_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_960_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_960_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_960_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_960_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_960_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_960_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_960_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_960_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_960_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_960_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_960_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_960_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_960_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_960_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_961_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_961_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_961_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_961_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_961_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_961_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_961_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_961_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_961_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_961_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_962_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_962_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_962_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_962_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_962_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_962_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_962_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_962_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_962_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_962_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_962_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_962_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_962_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_962_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_962_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_963_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_963_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_963_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_963_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_963_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_963_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_963_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_963_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_963_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_963_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_963_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_963_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_963_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_963_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_963_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_964_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_964_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_964_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_964_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_964_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_964_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_964_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_964_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_965_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_965_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_965_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_965_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_965_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_965_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_965_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_965_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_965_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_966_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_966_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_966_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_966_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_966_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_966_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_966_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_966_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_966_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_966_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_966_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_966_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_966_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_966_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_966_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_967_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_967_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_967_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_967_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_967_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_967_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_967_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_967_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_967_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_967_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_967_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_967_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_967_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_967_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_967_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_968_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_968_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_968_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_968_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_968_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_968_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_968_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_969_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_969_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_969_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_969_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_969_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_969_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_969_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_969_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_969_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_969_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_969_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_969_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_969_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_969_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_969_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_969_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_970_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_970_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_970_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_970_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_970_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_970_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_970_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_970_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_970_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_970_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_970_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_970_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_970_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_970_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_970_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_971_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_971_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_971_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_971_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_971_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_971_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_971_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_971_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_971_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_971_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_971_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_971_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_971_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_971_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_971_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_971_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_972_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_972_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_972_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_972_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_972_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_972_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_972_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_972_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_972_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_972_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_972_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_972_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_972_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_972_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_972_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_973_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_973_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_973_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_973_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_973_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_973_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_973_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_973_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_973_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_973_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_973_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_973_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_973_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_973_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_973_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_973_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_974_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_974_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_974_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_974_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_974_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_974_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_974_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_974_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_974_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_975_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_975_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_975_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_975_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_975_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_975_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_975_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_975_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_975_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_976_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_976_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_976_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_976_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_976_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_976_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_976_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_976_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_976_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_976_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_976_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_976_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_976_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_976_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_976_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_977_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_977_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_977_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_977_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_977_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_977_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_977_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_977_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_977_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_977_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_977_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_977_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_977_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_977_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_977_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_977_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_978_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_978_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_978_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_978_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_978_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_978_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_978_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_978_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_978_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_978_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_978_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_978_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_978_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_978_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_978_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_979_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_979_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_979_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_979_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_979_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_979_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_979_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_979_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_979_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_980_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_980_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_980_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_980_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_980_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_980_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_980_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_980_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_980_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_980_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_980_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_980_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_980_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_980_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_980_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_981_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_981_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_981_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_981_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_981_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_981_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_981_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_981_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_982_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_982_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_982_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_982_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_982_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_982_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_982_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_982_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_982_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_983_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_983_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_983_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_983_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_983_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_983_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_983_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_983_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_983_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_983_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_983_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_983_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_983_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_983_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_983_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_983_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_984_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_984_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_984_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_984_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_984_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_984_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_984_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_984_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_984_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_984_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_984_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_984_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_984_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_984_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_984_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_985_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_985_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_985_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_985_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_985_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_985_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_985_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_985_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_985_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_985_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_986_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_986_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_986_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_986_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_986_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_986_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_986_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_986_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_986_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_987_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_987_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_987_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_987_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_987_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_987_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_987_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_987_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_987_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_987_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_988_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_988_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_988_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_988_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_988_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_988_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_988_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_988_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_988_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_988_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_988_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_988_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_988_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_988_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_988_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_989_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_989_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_989_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_989_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_989_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_989_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_989_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_989_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_990_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_990_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_990_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_990_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_990_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_990_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_990_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_990_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_990_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_990_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_990_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_990_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_990_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_990_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_990_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_990_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_990_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_990_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_991_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_991_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_991_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_991_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_991_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_991_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_991_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_991_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_991_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_991_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_991_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_991_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_991_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_991_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_991_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_992_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_992_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_992_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_992_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_992_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_992_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_992_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_992_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_992_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_992_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_992_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_992_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_992_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_992_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_992_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_993_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_993_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_993_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_993_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_993_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_993_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_993_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_993_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_994_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_994_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_994_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_994_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_994_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_994_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_994_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_994_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_994_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_994_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_994_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_994_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_994_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_994_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_994_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_995_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_995_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_995_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_995_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_995_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_995_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_995_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_995_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_995_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_995_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_995_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_995_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_995_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_995_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_995_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_995_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_996_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_996_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_996_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_996_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_996_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_996_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_996_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_996_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_996_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_996_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_996_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_996_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_996_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_996_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_996_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_997_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_997_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_997_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_997_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_997_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_997_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_997_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_997_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_997_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_997_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_998_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_998_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_998_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_998_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_998_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_998_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_998_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_998_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_998_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_998_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_998_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_998_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_998_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_998_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_998_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_999_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_999_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_999_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_999_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_999_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_999_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_999_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_999_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_999_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_999_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_999_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_999_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_999_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_999_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_999_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_999_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_1000 ();
 sky130_fd_sc_hd__decap_3 PHY_1001 ();
 sky130_fd_sc_hd__decap_3 PHY_1002 ();
 sky130_fd_sc_hd__decap_3 PHY_1003 ();
 sky130_fd_sc_hd__decap_3 PHY_1004 ();
 sky130_fd_sc_hd__decap_3 PHY_1005 ();
 sky130_fd_sc_hd__decap_3 PHY_1006 ();
 sky130_fd_sc_hd__decap_3 PHY_1007 ();
 sky130_fd_sc_hd__decap_3 PHY_1008 ();
 sky130_fd_sc_hd__decap_3 PHY_1009 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_1010 ();
 sky130_fd_sc_hd__decap_3 PHY_1011 ();
 sky130_fd_sc_hd__decap_3 PHY_1012 ();
 sky130_fd_sc_hd__decap_3 PHY_1013 ();
 sky130_fd_sc_hd__decap_3 PHY_1014 ();
 sky130_fd_sc_hd__decap_3 PHY_1015 ();
 sky130_fd_sc_hd__decap_3 PHY_1016 ();
 sky130_fd_sc_hd__decap_3 PHY_1017 ();
 sky130_fd_sc_hd__decap_3 PHY_1018 ();
 sky130_fd_sc_hd__decap_3 PHY_1019 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_1020 ();
 sky130_fd_sc_hd__decap_3 PHY_1021 ();
 sky130_fd_sc_hd__decap_3 PHY_1022 ();
 sky130_fd_sc_hd__decap_3 PHY_1023 ();
 sky130_fd_sc_hd__decap_3 PHY_1024 ();
 sky130_fd_sc_hd__decap_3 PHY_1025 ();
 sky130_fd_sc_hd__decap_3 PHY_1026 ();
 sky130_fd_sc_hd__decap_3 PHY_1027 ();
 sky130_fd_sc_hd__decap_3 PHY_1028 ();
 sky130_fd_sc_hd__decap_3 PHY_1029 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_1030 ();
 sky130_fd_sc_hd__decap_3 PHY_1031 ();
 sky130_fd_sc_hd__decap_3 PHY_1032 ();
 sky130_fd_sc_hd__decap_3 PHY_1033 ();
 sky130_fd_sc_hd__decap_3 PHY_1034 ();
 sky130_fd_sc_hd__decap_3 PHY_1035 ();
 sky130_fd_sc_hd__decap_3 PHY_1036 ();
 sky130_fd_sc_hd__decap_3 PHY_1037 ();
 sky130_fd_sc_hd__decap_3 PHY_1038 ();
 sky130_fd_sc_hd__decap_3 PHY_1039 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_1040 ();
 sky130_fd_sc_hd__decap_3 PHY_1041 ();
 sky130_fd_sc_hd__decap_3 PHY_1042 ();
 sky130_fd_sc_hd__decap_3 PHY_1043 ();
 sky130_fd_sc_hd__decap_3 PHY_1044 ();
 sky130_fd_sc_hd__decap_3 PHY_1045 ();
 sky130_fd_sc_hd__decap_3 PHY_1046 ();
 sky130_fd_sc_hd__decap_3 PHY_1047 ();
 sky130_fd_sc_hd__decap_3 PHY_1048 ();
 sky130_fd_sc_hd__decap_3 PHY_1049 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_1050 ();
 sky130_fd_sc_hd__decap_3 PHY_1051 ();
 sky130_fd_sc_hd__decap_3 PHY_1052 ();
 sky130_fd_sc_hd__decap_3 PHY_1053 ();
 sky130_fd_sc_hd__decap_3 PHY_1054 ();
 sky130_fd_sc_hd__decap_3 PHY_1055 ();
 sky130_fd_sc_hd__decap_3 PHY_1056 ();
 sky130_fd_sc_hd__decap_3 PHY_1057 ();
 sky130_fd_sc_hd__decap_3 PHY_1058 ();
 sky130_fd_sc_hd__decap_3 PHY_1059 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_1060 ();
 sky130_fd_sc_hd__decap_3 PHY_1061 ();
 sky130_fd_sc_hd__decap_3 PHY_1062 ();
 sky130_fd_sc_hd__decap_3 PHY_1063 ();
 sky130_fd_sc_hd__decap_3 PHY_1064 ();
 sky130_fd_sc_hd__decap_3 PHY_1065 ();
 sky130_fd_sc_hd__decap_3 PHY_1066 ();
 sky130_fd_sc_hd__decap_3 PHY_1067 ();
 sky130_fd_sc_hd__decap_3 PHY_1068 ();
 sky130_fd_sc_hd__decap_3 PHY_1069 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_1070 ();
 sky130_fd_sc_hd__decap_3 PHY_1071 ();
 sky130_fd_sc_hd__decap_3 PHY_1072 ();
 sky130_fd_sc_hd__decap_3 PHY_1073 ();
 sky130_fd_sc_hd__decap_3 PHY_1074 ();
 sky130_fd_sc_hd__decap_3 PHY_1075 ();
 sky130_fd_sc_hd__decap_3 PHY_1076 ();
 sky130_fd_sc_hd__decap_3 PHY_1077 ();
 sky130_fd_sc_hd__decap_3 PHY_1078 ();
 sky130_fd_sc_hd__decap_3 PHY_1079 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_1080 ();
 sky130_fd_sc_hd__decap_3 PHY_1081 ();
 sky130_fd_sc_hd__decap_3 PHY_1082 ();
 sky130_fd_sc_hd__decap_3 PHY_1083 ();
 sky130_fd_sc_hd__decap_3 PHY_1084 ();
 sky130_fd_sc_hd__decap_3 PHY_1085 ();
 sky130_fd_sc_hd__decap_3 PHY_1086 ();
 sky130_fd_sc_hd__decap_3 PHY_1087 ();
 sky130_fd_sc_hd__decap_3 PHY_1088 ();
 sky130_fd_sc_hd__decap_3 PHY_1089 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_1090 ();
 sky130_fd_sc_hd__decap_3 PHY_1091 ();
 sky130_fd_sc_hd__decap_3 PHY_1092 ();
 sky130_fd_sc_hd__decap_3 PHY_1093 ();
 sky130_fd_sc_hd__decap_3 PHY_1094 ();
 sky130_fd_sc_hd__decap_3 PHY_1095 ();
 sky130_fd_sc_hd__decap_3 PHY_1096 ();
 sky130_fd_sc_hd__decap_3 PHY_1097 ();
 sky130_fd_sc_hd__decap_3 PHY_1098 ();
 sky130_fd_sc_hd__decap_3 PHY_1099 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_1100 ();
 sky130_fd_sc_hd__decap_3 PHY_1101 ();
 sky130_fd_sc_hd__decap_3 PHY_1102 ();
 sky130_fd_sc_hd__decap_3 PHY_1103 ();
 sky130_fd_sc_hd__decap_3 PHY_1104 ();
 sky130_fd_sc_hd__decap_3 PHY_1105 ();
 sky130_fd_sc_hd__decap_3 PHY_1106 ();
 sky130_fd_sc_hd__decap_3 PHY_1107 ();
 sky130_fd_sc_hd__decap_3 PHY_1108 ();
 sky130_fd_sc_hd__decap_3 PHY_1109 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_1110 ();
 sky130_fd_sc_hd__decap_3 PHY_1111 ();
 sky130_fd_sc_hd__decap_3 PHY_1112 ();
 sky130_fd_sc_hd__decap_3 PHY_1113 ();
 sky130_fd_sc_hd__decap_3 PHY_1114 ();
 sky130_fd_sc_hd__decap_3 PHY_1115 ();
 sky130_fd_sc_hd__decap_3 PHY_1116 ();
 sky130_fd_sc_hd__decap_3 PHY_1117 ();
 sky130_fd_sc_hd__decap_3 PHY_1118 ();
 sky130_fd_sc_hd__decap_3 PHY_1119 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_1120 ();
 sky130_fd_sc_hd__decap_3 PHY_1121 ();
 sky130_fd_sc_hd__decap_3 PHY_1122 ();
 sky130_fd_sc_hd__decap_3 PHY_1123 ();
 sky130_fd_sc_hd__decap_3 PHY_1124 ();
 sky130_fd_sc_hd__decap_3 PHY_1125 ();
 sky130_fd_sc_hd__decap_3 PHY_1126 ();
 sky130_fd_sc_hd__decap_3 PHY_1127 ();
 sky130_fd_sc_hd__decap_3 PHY_1128 ();
 sky130_fd_sc_hd__decap_3 PHY_1129 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_1130 ();
 sky130_fd_sc_hd__decap_3 PHY_1131 ();
 sky130_fd_sc_hd__decap_3 PHY_1132 ();
 sky130_fd_sc_hd__decap_3 PHY_1133 ();
 sky130_fd_sc_hd__decap_3 PHY_1134 ();
 sky130_fd_sc_hd__decap_3 PHY_1135 ();
 sky130_fd_sc_hd__decap_3 PHY_1136 ();
 sky130_fd_sc_hd__decap_3 PHY_1137 ();
 sky130_fd_sc_hd__decap_3 PHY_1138 ();
 sky130_fd_sc_hd__decap_3 PHY_1139 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_1140 ();
 sky130_fd_sc_hd__decap_3 PHY_1141 ();
 sky130_fd_sc_hd__decap_3 PHY_1142 ();
 sky130_fd_sc_hd__decap_3 PHY_1143 ();
 sky130_fd_sc_hd__decap_3 PHY_1144 ();
 sky130_fd_sc_hd__decap_3 PHY_1145 ();
 sky130_fd_sc_hd__decap_3 PHY_1146 ();
 sky130_fd_sc_hd__decap_3 PHY_1147 ();
 sky130_fd_sc_hd__decap_3 PHY_1148 ();
 sky130_fd_sc_hd__decap_3 PHY_1149 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_1150 ();
 sky130_fd_sc_hd__decap_3 PHY_1151 ();
 sky130_fd_sc_hd__decap_3 PHY_1152 ();
 sky130_fd_sc_hd__decap_3 PHY_1153 ();
 sky130_fd_sc_hd__decap_3 PHY_1154 ();
 sky130_fd_sc_hd__decap_3 PHY_1155 ();
 sky130_fd_sc_hd__decap_3 PHY_1156 ();
 sky130_fd_sc_hd__decap_3 PHY_1157 ();
 sky130_fd_sc_hd__decap_3 PHY_1158 ();
 sky130_fd_sc_hd__decap_3 PHY_1159 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_1160 ();
 sky130_fd_sc_hd__decap_3 PHY_1161 ();
 sky130_fd_sc_hd__decap_3 PHY_1162 ();
 sky130_fd_sc_hd__decap_3 PHY_1163 ();
 sky130_fd_sc_hd__decap_3 PHY_1164 ();
 sky130_fd_sc_hd__decap_3 PHY_1165 ();
 sky130_fd_sc_hd__decap_3 PHY_1166 ();
 sky130_fd_sc_hd__decap_3 PHY_1167 ();
 sky130_fd_sc_hd__decap_3 PHY_1168 ();
 sky130_fd_sc_hd__decap_3 PHY_1169 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_1170 ();
 sky130_fd_sc_hd__decap_3 PHY_1171 ();
 sky130_fd_sc_hd__decap_3 PHY_1172 ();
 sky130_fd_sc_hd__decap_3 PHY_1173 ();
 sky130_fd_sc_hd__decap_3 PHY_1174 ();
 sky130_fd_sc_hd__decap_3 PHY_1175 ();
 sky130_fd_sc_hd__decap_3 PHY_1176 ();
 sky130_fd_sc_hd__decap_3 PHY_1177 ();
 sky130_fd_sc_hd__decap_3 PHY_1178 ();
 sky130_fd_sc_hd__decap_3 PHY_1179 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_1180 ();
 sky130_fd_sc_hd__decap_3 PHY_1181 ();
 sky130_fd_sc_hd__decap_3 PHY_1182 ();
 sky130_fd_sc_hd__decap_3 PHY_1183 ();
 sky130_fd_sc_hd__decap_3 PHY_1184 ();
 sky130_fd_sc_hd__decap_3 PHY_1185 ();
 sky130_fd_sc_hd__decap_3 PHY_1186 ();
 sky130_fd_sc_hd__decap_3 PHY_1187 ();
 sky130_fd_sc_hd__decap_3 PHY_1188 ();
 sky130_fd_sc_hd__decap_3 PHY_1189 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_1190 ();
 sky130_fd_sc_hd__decap_3 PHY_1191 ();
 sky130_fd_sc_hd__decap_3 PHY_1192 ();
 sky130_fd_sc_hd__decap_3 PHY_1193 ();
 sky130_fd_sc_hd__decap_3 PHY_1194 ();
 sky130_fd_sc_hd__decap_3 PHY_1195 ();
 sky130_fd_sc_hd__decap_3 PHY_1196 ();
 sky130_fd_sc_hd__decap_3 PHY_1197 ();
 sky130_fd_sc_hd__decap_3 PHY_1198 ();
 sky130_fd_sc_hd__decap_3 PHY_1199 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_1200 ();
 sky130_fd_sc_hd__decap_3 PHY_1201 ();
 sky130_fd_sc_hd__decap_3 PHY_1202 ();
 sky130_fd_sc_hd__decap_3 PHY_1203 ();
 sky130_fd_sc_hd__decap_3 PHY_1204 ();
 sky130_fd_sc_hd__decap_3 PHY_1205 ();
 sky130_fd_sc_hd__decap_3 PHY_1206 ();
 sky130_fd_sc_hd__decap_3 PHY_1207 ();
 sky130_fd_sc_hd__decap_3 PHY_1208 ();
 sky130_fd_sc_hd__decap_3 PHY_1209 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_1210 ();
 sky130_fd_sc_hd__decap_3 PHY_1211 ();
 sky130_fd_sc_hd__decap_3 PHY_1212 ();
 sky130_fd_sc_hd__decap_3 PHY_1213 ();
 sky130_fd_sc_hd__decap_3 PHY_1214 ();
 sky130_fd_sc_hd__decap_3 PHY_1215 ();
 sky130_fd_sc_hd__decap_3 PHY_1216 ();
 sky130_fd_sc_hd__decap_3 PHY_1217 ();
 sky130_fd_sc_hd__decap_3 PHY_1218 ();
 sky130_fd_sc_hd__decap_3 PHY_1219 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_1220 ();
 sky130_fd_sc_hd__decap_3 PHY_1221 ();
 sky130_fd_sc_hd__decap_3 PHY_1222 ();
 sky130_fd_sc_hd__decap_3 PHY_1223 ();
 sky130_fd_sc_hd__decap_3 PHY_1224 ();
 sky130_fd_sc_hd__decap_3 PHY_1225 ();
 sky130_fd_sc_hd__decap_3 PHY_1226 ();
 sky130_fd_sc_hd__decap_3 PHY_1227 ();
 sky130_fd_sc_hd__decap_3 PHY_1228 ();
 sky130_fd_sc_hd__decap_3 PHY_1229 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_1230 ();
 sky130_fd_sc_hd__decap_3 PHY_1231 ();
 sky130_fd_sc_hd__decap_3 PHY_1232 ();
 sky130_fd_sc_hd__decap_3 PHY_1233 ();
 sky130_fd_sc_hd__decap_3 PHY_1234 ();
 sky130_fd_sc_hd__decap_3 PHY_1235 ();
 sky130_fd_sc_hd__decap_3 PHY_1236 ();
 sky130_fd_sc_hd__decap_3 PHY_1237 ();
 sky130_fd_sc_hd__decap_3 PHY_1238 ();
 sky130_fd_sc_hd__decap_3 PHY_1239 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_1240 ();
 sky130_fd_sc_hd__decap_3 PHY_1241 ();
 sky130_fd_sc_hd__decap_3 PHY_1242 ();
 sky130_fd_sc_hd__decap_3 PHY_1243 ();
 sky130_fd_sc_hd__decap_3 PHY_1244 ();
 sky130_fd_sc_hd__decap_3 PHY_1245 ();
 sky130_fd_sc_hd__decap_3 PHY_1246 ();
 sky130_fd_sc_hd__decap_3 PHY_1247 ();
 sky130_fd_sc_hd__decap_3 PHY_1248 ();
 sky130_fd_sc_hd__decap_3 PHY_1249 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_1250 ();
 sky130_fd_sc_hd__decap_3 PHY_1251 ();
 sky130_fd_sc_hd__decap_3 PHY_1252 ();
 sky130_fd_sc_hd__decap_3 PHY_1253 ();
 sky130_fd_sc_hd__decap_3 PHY_1254 ();
 sky130_fd_sc_hd__decap_3 PHY_1255 ();
 sky130_fd_sc_hd__decap_3 PHY_1256 ();
 sky130_fd_sc_hd__decap_3 PHY_1257 ();
 sky130_fd_sc_hd__decap_3 PHY_1258 ();
 sky130_fd_sc_hd__decap_3 PHY_1259 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_1260 ();
 sky130_fd_sc_hd__decap_3 PHY_1261 ();
 sky130_fd_sc_hd__decap_3 PHY_1262 ();
 sky130_fd_sc_hd__decap_3 PHY_1263 ();
 sky130_fd_sc_hd__decap_3 PHY_1264 ();
 sky130_fd_sc_hd__decap_3 PHY_1265 ();
 sky130_fd_sc_hd__decap_3 PHY_1266 ();
 sky130_fd_sc_hd__decap_3 PHY_1267 ();
 sky130_fd_sc_hd__decap_3 PHY_1268 ();
 sky130_fd_sc_hd__decap_3 PHY_1269 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_1270 ();
 sky130_fd_sc_hd__decap_3 PHY_1271 ();
 sky130_fd_sc_hd__decap_3 PHY_1272 ();
 sky130_fd_sc_hd__decap_3 PHY_1273 ();
 sky130_fd_sc_hd__decap_3 PHY_1274 ();
 sky130_fd_sc_hd__decap_3 PHY_1275 ();
 sky130_fd_sc_hd__decap_3 PHY_1276 ();
 sky130_fd_sc_hd__decap_3 PHY_1277 ();
 sky130_fd_sc_hd__decap_3 PHY_1278 ();
 sky130_fd_sc_hd__decap_3 PHY_1279 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_1280 ();
 sky130_fd_sc_hd__decap_3 PHY_1281 ();
 sky130_fd_sc_hd__decap_3 PHY_1282 ();
 sky130_fd_sc_hd__decap_3 PHY_1283 ();
 sky130_fd_sc_hd__decap_3 PHY_1284 ();
 sky130_fd_sc_hd__decap_3 PHY_1285 ();
 sky130_fd_sc_hd__decap_3 PHY_1286 ();
 sky130_fd_sc_hd__decap_3 PHY_1287 ();
 sky130_fd_sc_hd__decap_3 PHY_1288 ();
 sky130_fd_sc_hd__decap_3 PHY_1289 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_1290 ();
 sky130_fd_sc_hd__decap_3 PHY_1291 ();
 sky130_fd_sc_hd__decap_3 PHY_1292 ();
 sky130_fd_sc_hd__decap_3 PHY_1293 ();
 sky130_fd_sc_hd__decap_3 PHY_1294 ();
 sky130_fd_sc_hd__decap_3 PHY_1295 ();
 sky130_fd_sc_hd__decap_3 PHY_1296 ();
 sky130_fd_sc_hd__decap_3 PHY_1297 ();
 sky130_fd_sc_hd__decap_3 PHY_1298 ();
 sky130_fd_sc_hd__decap_3 PHY_1299 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_1300 ();
 sky130_fd_sc_hd__decap_3 PHY_1301 ();
 sky130_fd_sc_hd__decap_3 PHY_1302 ();
 sky130_fd_sc_hd__decap_3 PHY_1303 ();
 sky130_fd_sc_hd__decap_3 PHY_1304 ();
 sky130_fd_sc_hd__decap_3 PHY_1305 ();
 sky130_fd_sc_hd__decap_3 PHY_1306 ();
 sky130_fd_sc_hd__decap_3 PHY_1307 ();
 sky130_fd_sc_hd__decap_3 PHY_1308 ();
 sky130_fd_sc_hd__decap_3 PHY_1309 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_1310 ();
 sky130_fd_sc_hd__decap_3 PHY_1311 ();
 sky130_fd_sc_hd__decap_3 PHY_1312 ();
 sky130_fd_sc_hd__decap_3 PHY_1313 ();
 sky130_fd_sc_hd__decap_3 PHY_1314 ();
 sky130_fd_sc_hd__decap_3 PHY_1315 ();
 sky130_fd_sc_hd__decap_3 PHY_1316 ();
 sky130_fd_sc_hd__decap_3 PHY_1317 ();
 sky130_fd_sc_hd__decap_3 PHY_1318 ();
 sky130_fd_sc_hd__decap_3 PHY_1319 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_1320 ();
 sky130_fd_sc_hd__decap_3 PHY_1321 ();
 sky130_fd_sc_hd__decap_3 PHY_1322 ();
 sky130_fd_sc_hd__decap_3 PHY_1323 ();
 sky130_fd_sc_hd__decap_3 PHY_1324 ();
 sky130_fd_sc_hd__decap_3 PHY_1325 ();
 sky130_fd_sc_hd__decap_3 PHY_1326 ();
 sky130_fd_sc_hd__decap_3 PHY_1327 ();
 sky130_fd_sc_hd__decap_3 PHY_1328 ();
 sky130_fd_sc_hd__decap_3 PHY_1329 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_1330 ();
 sky130_fd_sc_hd__decap_3 PHY_1331 ();
 sky130_fd_sc_hd__decap_3 PHY_1332 ();
 sky130_fd_sc_hd__decap_3 PHY_1333 ();
 sky130_fd_sc_hd__decap_3 PHY_1334 ();
 sky130_fd_sc_hd__decap_3 PHY_1335 ();
 sky130_fd_sc_hd__decap_3 PHY_1336 ();
 sky130_fd_sc_hd__decap_3 PHY_1337 ();
 sky130_fd_sc_hd__decap_3 PHY_1338 ();
 sky130_fd_sc_hd__decap_3 PHY_1339 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_1340 ();
 sky130_fd_sc_hd__decap_3 PHY_1341 ();
 sky130_fd_sc_hd__decap_3 PHY_1342 ();
 sky130_fd_sc_hd__decap_3 PHY_1343 ();
 sky130_fd_sc_hd__decap_3 PHY_1344 ();
 sky130_fd_sc_hd__decap_3 PHY_1345 ();
 sky130_fd_sc_hd__decap_3 PHY_1346 ();
 sky130_fd_sc_hd__decap_3 PHY_1347 ();
 sky130_fd_sc_hd__decap_3 PHY_1348 ();
 sky130_fd_sc_hd__decap_3 PHY_1349 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_1350 ();
 sky130_fd_sc_hd__decap_3 PHY_1351 ();
 sky130_fd_sc_hd__decap_3 PHY_1352 ();
 sky130_fd_sc_hd__decap_3 PHY_1353 ();
 sky130_fd_sc_hd__decap_3 PHY_1354 ();
 sky130_fd_sc_hd__decap_3 PHY_1355 ();
 sky130_fd_sc_hd__decap_3 PHY_1356 ();
 sky130_fd_sc_hd__decap_3 PHY_1357 ();
 sky130_fd_sc_hd__decap_3 PHY_1358 ();
 sky130_fd_sc_hd__decap_3 PHY_1359 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_1360 ();
 sky130_fd_sc_hd__decap_3 PHY_1361 ();
 sky130_fd_sc_hd__decap_3 PHY_1362 ();
 sky130_fd_sc_hd__decap_3 PHY_1363 ();
 sky130_fd_sc_hd__decap_3 PHY_1364 ();
 sky130_fd_sc_hd__decap_3 PHY_1365 ();
 sky130_fd_sc_hd__decap_3 PHY_1366 ();
 sky130_fd_sc_hd__decap_3 PHY_1367 ();
 sky130_fd_sc_hd__decap_3 PHY_1368 ();
 sky130_fd_sc_hd__decap_3 PHY_1369 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_1370 ();
 sky130_fd_sc_hd__decap_3 PHY_1371 ();
 sky130_fd_sc_hd__decap_3 PHY_1372 ();
 sky130_fd_sc_hd__decap_3 PHY_1373 ();
 sky130_fd_sc_hd__decap_3 PHY_1374 ();
 sky130_fd_sc_hd__decap_3 PHY_1375 ();
 sky130_fd_sc_hd__decap_3 PHY_1376 ();
 sky130_fd_sc_hd__decap_3 PHY_1377 ();
 sky130_fd_sc_hd__decap_3 PHY_1378 ();
 sky130_fd_sc_hd__decap_3 PHY_1379 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_1380 ();
 sky130_fd_sc_hd__decap_3 PHY_1381 ();
 sky130_fd_sc_hd__decap_3 PHY_1382 ();
 sky130_fd_sc_hd__decap_3 PHY_1383 ();
 sky130_fd_sc_hd__decap_3 PHY_1384 ();
 sky130_fd_sc_hd__decap_3 PHY_1385 ();
 sky130_fd_sc_hd__decap_3 PHY_1386 ();
 sky130_fd_sc_hd__decap_3 PHY_1387 ();
 sky130_fd_sc_hd__decap_3 PHY_1388 ();
 sky130_fd_sc_hd__decap_3 PHY_1389 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_1390 ();
 sky130_fd_sc_hd__decap_3 PHY_1391 ();
 sky130_fd_sc_hd__decap_3 PHY_1392 ();
 sky130_fd_sc_hd__decap_3 PHY_1393 ();
 sky130_fd_sc_hd__decap_3 PHY_1394 ();
 sky130_fd_sc_hd__decap_3 PHY_1395 ();
 sky130_fd_sc_hd__decap_3 PHY_1396 ();
 sky130_fd_sc_hd__decap_3 PHY_1397 ();
 sky130_fd_sc_hd__decap_3 PHY_1398 ();
 sky130_fd_sc_hd__decap_3 PHY_1399 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_1400 ();
 sky130_fd_sc_hd__decap_3 PHY_1401 ();
 sky130_fd_sc_hd__decap_3 PHY_1402 ();
 sky130_fd_sc_hd__decap_3 PHY_1403 ();
 sky130_fd_sc_hd__decap_3 PHY_1404 ();
 sky130_fd_sc_hd__decap_3 PHY_1405 ();
 sky130_fd_sc_hd__decap_3 PHY_1406 ();
 sky130_fd_sc_hd__decap_3 PHY_1407 ();
 sky130_fd_sc_hd__decap_3 PHY_1408 ();
 sky130_fd_sc_hd__decap_3 PHY_1409 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_1410 ();
 sky130_fd_sc_hd__decap_3 PHY_1411 ();
 sky130_fd_sc_hd__decap_3 PHY_1412 ();
 sky130_fd_sc_hd__decap_3 PHY_1413 ();
 sky130_fd_sc_hd__decap_3 PHY_1414 ();
 sky130_fd_sc_hd__decap_3 PHY_1415 ();
 sky130_fd_sc_hd__decap_3 PHY_1416 ();
 sky130_fd_sc_hd__decap_3 PHY_1417 ();
 sky130_fd_sc_hd__decap_3 PHY_1418 ();
 sky130_fd_sc_hd__decap_3 PHY_1419 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_1420 ();
 sky130_fd_sc_hd__decap_3 PHY_1421 ();
 sky130_fd_sc_hd__decap_3 PHY_1422 ();
 sky130_fd_sc_hd__decap_3 PHY_1423 ();
 sky130_fd_sc_hd__decap_3 PHY_1424 ();
 sky130_fd_sc_hd__decap_3 PHY_1425 ();
 sky130_fd_sc_hd__decap_3 PHY_1426 ();
 sky130_fd_sc_hd__decap_3 PHY_1427 ();
 sky130_fd_sc_hd__decap_3 PHY_1428 ();
 sky130_fd_sc_hd__decap_3 PHY_1429 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_1430 ();
 sky130_fd_sc_hd__decap_3 PHY_1431 ();
 sky130_fd_sc_hd__decap_3 PHY_1432 ();
 sky130_fd_sc_hd__decap_3 PHY_1433 ();
 sky130_fd_sc_hd__decap_3 PHY_1434 ();
 sky130_fd_sc_hd__decap_3 PHY_1435 ();
 sky130_fd_sc_hd__decap_3 PHY_1436 ();
 sky130_fd_sc_hd__decap_3 PHY_1437 ();
 sky130_fd_sc_hd__decap_3 PHY_1438 ();
 sky130_fd_sc_hd__decap_3 PHY_1439 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_1440 ();
 sky130_fd_sc_hd__decap_3 PHY_1441 ();
 sky130_fd_sc_hd__decap_3 PHY_1442 ();
 sky130_fd_sc_hd__decap_3 PHY_1443 ();
 sky130_fd_sc_hd__decap_3 PHY_1444 ();
 sky130_fd_sc_hd__decap_3 PHY_1445 ();
 sky130_fd_sc_hd__decap_3 PHY_1446 ();
 sky130_fd_sc_hd__decap_3 PHY_1447 ();
 sky130_fd_sc_hd__decap_3 PHY_1448 ();
 sky130_fd_sc_hd__decap_3 PHY_1449 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_1450 ();
 sky130_fd_sc_hd__decap_3 PHY_1451 ();
 sky130_fd_sc_hd__decap_3 PHY_1452 ();
 sky130_fd_sc_hd__decap_3 PHY_1453 ();
 sky130_fd_sc_hd__decap_3 PHY_1454 ();
 sky130_fd_sc_hd__decap_3 PHY_1455 ();
 sky130_fd_sc_hd__decap_3 PHY_1456 ();
 sky130_fd_sc_hd__decap_3 PHY_1457 ();
 sky130_fd_sc_hd__decap_3 PHY_1458 ();
 sky130_fd_sc_hd__decap_3 PHY_1459 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_1460 ();
 sky130_fd_sc_hd__decap_3 PHY_1461 ();
 sky130_fd_sc_hd__decap_3 PHY_1462 ();
 sky130_fd_sc_hd__decap_3 PHY_1463 ();
 sky130_fd_sc_hd__decap_3 PHY_1464 ();
 sky130_fd_sc_hd__decap_3 PHY_1465 ();
 sky130_fd_sc_hd__decap_3 PHY_1466 ();
 sky130_fd_sc_hd__decap_3 PHY_1467 ();
 sky130_fd_sc_hd__decap_3 PHY_1468 ();
 sky130_fd_sc_hd__decap_3 PHY_1469 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_1470 ();
 sky130_fd_sc_hd__decap_3 PHY_1471 ();
 sky130_fd_sc_hd__decap_3 PHY_1472 ();
 sky130_fd_sc_hd__decap_3 PHY_1473 ();
 sky130_fd_sc_hd__decap_3 PHY_1474 ();
 sky130_fd_sc_hd__decap_3 PHY_1475 ();
 sky130_fd_sc_hd__decap_3 PHY_1476 ();
 sky130_fd_sc_hd__decap_3 PHY_1477 ();
 sky130_fd_sc_hd__decap_3 PHY_1478 ();
 sky130_fd_sc_hd__decap_3 PHY_1479 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_1480 ();
 sky130_fd_sc_hd__decap_3 PHY_1481 ();
 sky130_fd_sc_hd__decap_3 PHY_1482 ();
 sky130_fd_sc_hd__decap_3 PHY_1483 ();
 sky130_fd_sc_hd__decap_3 PHY_1484 ();
 sky130_fd_sc_hd__decap_3 PHY_1485 ();
 sky130_fd_sc_hd__decap_3 PHY_1486 ();
 sky130_fd_sc_hd__decap_3 PHY_1487 ();
 sky130_fd_sc_hd__decap_3 PHY_1488 ();
 sky130_fd_sc_hd__decap_3 PHY_1489 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_1490 ();
 sky130_fd_sc_hd__decap_3 PHY_1491 ();
 sky130_fd_sc_hd__decap_3 PHY_1492 ();
 sky130_fd_sc_hd__decap_3 PHY_1493 ();
 sky130_fd_sc_hd__decap_3 PHY_1494 ();
 sky130_fd_sc_hd__decap_3 PHY_1495 ();
 sky130_fd_sc_hd__decap_3 PHY_1496 ();
 sky130_fd_sc_hd__decap_3 PHY_1497 ();
 sky130_fd_sc_hd__decap_3 PHY_1498 ();
 sky130_fd_sc_hd__decap_3 PHY_1499 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_1500 ();
 sky130_fd_sc_hd__decap_3 PHY_1501 ();
 sky130_fd_sc_hd__decap_3 PHY_1502 ();
 sky130_fd_sc_hd__decap_3 PHY_1503 ();
 sky130_fd_sc_hd__decap_3 PHY_1504 ();
 sky130_fd_sc_hd__decap_3 PHY_1505 ();
 sky130_fd_sc_hd__decap_3 PHY_1506 ();
 sky130_fd_sc_hd__decap_3 PHY_1507 ();
 sky130_fd_sc_hd__decap_3 PHY_1508 ();
 sky130_fd_sc_hd__decap_3 PHY_1509 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_1510 ();
 sky130_fd_sc_hd__decap_3 PHY_1511 ();
 sky130_fd_sc_hd__decap_3 PHY_1512 ();
 sky130_fd_sc_hd__decap_3 PHY_1513 ();
 sky130_fd_sc_hd__decap_3 PHY_1514 ();
 sky130_fd_sc_hd__decap_3 PHY_1515 ();
 sky130_fd_sc_hd__decap_3 PHY_1516 ();
 sky130_fd_sc_hd__decap_3 PHY_1517 ();
 sky130_fd_sc_hd__decap_3 PHY_1518 ();
 sky130_fd_sc_hd__decap_3 PHY_1519 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_1520 ();
 sky130_fd_sc_hd__decap_3 PHY_1521 ();
 sky130_fd_sc_hd__decap_3 PHY_1522 ();
 sky130_fd_sc_hd__decap_3 PHY_1523 ();
 sky130_fd_sc_hd__decap_3 PHY_1524 ();
 sky130_fd_sc_hd__decap_3 PHY_1525 ();
 sky130_fd_sc_hd__decap_3 PHY_1526 ();
 sky130_fd_sc_hd__decap_3 PHY_1527 ();
 sky130_fd_sc_hd__decap_3 PHY_1528 ();
 sky130_fd_sc_hd__decap_3 PHY_1529 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_1530 ();
 sky130_fd_sc_hd__decap_3 PHY_1531 ();
 sky130_fd_sc_hd__decap_3 PHY_1532 ();
 sky130_fd_sc_hd__decap_3 PHY_1533 ();
 sky130_fd_sc_hd__decap_3 PHY_1534 ();
 sky130_fd_sc_hd__decap_3 PHY_1535 ();
 sky130_fd_sc_hd__decap_3 PHY_1536 ();
 sky130_fd_sc_hd__decap_3 PHY_1537 ();
 sky130_fd_sc_hd__decap_3 PHY_1538 ();
 sky130_fd_sc_hd__decap_3 PHY_1539 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_1540 ();
 sky130_fd_sc_hd__decap_3 PHY_1541 ();
 sky130_fd_sc_hd__decap_3 PHY_1542 ();
 sky130_fd_sc_hd__decap_3 PHY_1543 ();
 sky130_fd_sc_hd__decap_3 PHY_1544 ();
 sky130_fd_sc_hd__decap_3 PHY_1545 ();
 sky130_fd_sc_hd__decap_3 PHY_1546 ();
 sky130_fd_sc_hd__decap_3 PHY_1547 ();
 sky130_fd_sc_hd__decap_3 PHY_1548 ();
 sky130_fd_sc_hd__decap_3 PHY_1549 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_1550 ();
 sky130_fd_sc_hd__decap_3 PHY_1551 ();
 sky130_fd_sc_hd__decap_3 PHY_1552 ();
 sky130_fd_sc_hd__decap_3 PHY_1553 ();
 sky130_fd_sc_hd__decap_3 PHY_1554 ();
 sky130_fd_sc_hd__decap_3 PHY_1555 ();
 sky130_fd_sc_hd__decap_3 PHY_1556 ();
 sky130_fd_sc_hd__decap_3 PHY_1557 ();
 sky130_fd_sc_hd__decap_3 PHY_1558 ();
 sky130_fd_sc_hd__decap_3 PHY_1559 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_1560 ();
 sky130_fd_sc_hd__decap_3 PHY_1561 ();
 sky130_fd_sc_hd__decap_3 PHY_1562 ();
 sky130_fd_sc_hd__decap_3 PHY_1563 ();
 sky130_fd_sc_hd__decap_3 PHY_1564 ();
 sky130_fd_sc_hd__decap_3 PHY_1565 ();
 sky130_fd_sc_hd__decap_3 PHY_1566 ();
 sky130_fd_sc_hd__decap_3 PHY_1567 ();
 sky130_fd_sc_hd__decap_3 PHY_1568 ();
 sky130_fd_sc_hd__decap_3 PHY_1569 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_1570 ();
 sky130_fd_sc_hd__decap_3 PHY_1571 ();
 sky130_fd_sc_hd__decap_3 PHY_1572 ();
 sky130_fd_sc_hd__decap_3 PHY_1573 ();
 sky130_fd_sc_hd__decap_3 PHY_1574 ();
 sky130_fd_sc_hd__decap_3 PHY_1575 ();
 sky130_fd_sc_hd__decap_3 PHY_1576 ();
 sky130_fd_sc_hd__decap_3 PHY_1577 ();
 sky130_fd_sc_hd__decap_3 PHY_1578 ();
 sky130_fd_sc_hd__decap_3 PHY_1579 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_1580 ();
 sky130_fd_sc_hd__decap_3 PHY_1581 ();
 sky130_fd_sc_hd__decap_3 PHY_1582 ();
 sky130_fd_sc_hd__decap_3 PHY_1583 ();
 sky130_fd_sc_hd__decap_3 PHY_1584 ();
 sky130_fd_sc_hd__decap_3 PHY_1585 ();
 sky130_fd_sc_hd__decap_3 PHY_1586 ();
 sky130_fd_sc_hd__decap_3 PHY_1587 ();
 sky130_fd_sc_hd__decap_3 PHY_1588 ();
 sky130_fd_sc_hd__decap_3 PHY_1589 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_1590 ();
 sky130_fd_sc_hd__decap_3 PHY_1591 ();
 sky130_fd_sc_hd__decap_3 PHY_1592 ();
 sky130_fd_sc_hd__decap_3 PHY_1593 ();
 sky130_fd_sc_hd__decap_3 PHY_1594 ();
 sky130_fd_sc_hd__decap_3 PHY_1595 ();
 sky130_fd_sc_hd__decap_3 PHY_1596 ();
 sky130_fd_sc_hd__decap_3 PHY_1597 ();
 sky130_fd_sc_hd__decap_3 PHY_1598 ();
 sky130_fd_sc_hd__decap_3 PHY_1599 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_1600 ();
 sky130_fd_sc_hd__decap_3 PHY_1601 ();
 sky130_fd_sc_hd__decap_3 PHY_1602 ();
 sky130_fd_sc_hd__decap_3 PHY_1603 ();
 sky130_fd_sc_hd__decap_3 PHY_1604 ();
 sky130_fd_sc_hd__decap_3 PHY_1605 ();
 sky130_fd_sc_hd__decap_3 PHY_1606 ();
 sky130_fd_sc_hd__decap_3 PHY_1607 ();
 sky130_fd_sc_hd__decap_3 PHY_1608 ();
 sky130_fd_sc_hd__decap_3 PHY_1609 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_1610 ();
 sky130_fd_sc_hd__decap_3 PHY_1611 ();
 sky130_fd_sc_hd__decap_3 PHY_1612 ();
 sky130_fd_sc_hd__decap_3 PHY_1613 ();
 sky130_fd_sc_hd__decap_3 PHY_1614 ();
 sky130_fd_sc_hd__decap_3 PHY_1615 ();
 sky130_fd_sc_hd__decap_3 PHY_1616 ();
 sky130_fd_sc_hd__decap_3 PHY_1617 ();
 sky130_fd_sc_hd__decap_3 PHY_1618 ();
 sky130_fd_sc_hd__decap_3 PHY_1619 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_1620 ();
 sky130_fd_sc_hd__decap_3 PHY_1621 ();
 sky130_fd_sc_hd__decap_3 PHY_1622 ();
 sky130_fd_sc_hd__decap_3 PHY_1623 ();
 sky130_fd_sc_hd__decap_3 PHY_1624 ();
 sky130_fd_sc_hd__decap_3 PHY_1625 ();
 sky130_fd_sc_hd__decap_3 PHY_1626 ();
 sky130_fd_sc_hd__decap_3 PHY_1627 ();
 sky130_fd_sc_hd__decap_3 PHY_1628 ();
 sky130_fd_sc_hd__decap_3 PHY_1629 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_1630 ();
 sky130_fd_sc_hd__decap_3 PHY_1631 ();
 sky130_fd_sc_hd__decap_3 PHY_1632 ();
 sky130_fd_sc_hd__decap_3 PHY_1633 ();
 sky130_fd_sc_hd__decap_3 PHY_1634 ();
 sky130_fd_sc_hd__decap_3 PHY_1635 ();
 sky130_fd_sc_hd__decap_3 PHY_1636 ();
 sky130_fd_sc_hd__decap_3 PHY_1637 ();
 sky130_fd_sc_hd__decap_3 PHY_1638 ();
 sky130_fd_sc_hd__decap_3 PHY_1639 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_1640 ();
 sky130_fd_sc_hd__decap_3 PHY_1641 ();
 sky130_fd_sc_hd__decap_3 PHY_1642 ();
 sky130_fd_sc_hd__decap_3 PHY_1643 ();
 sky130_fd_sc_hd__decap_3 PHY_1644 ();
 sky130_fd_sc_hd__decap_3 PHY_1645 ();
 sky130_fd_sc_hd__decap_3 PHY_1646 ();
 sky130_fd_sc_hd__decap_3 PHY_1647 ();
 sky130_fd_sc_hd__decap_3 PHY_1648 ();
 sky130_fd_sc_hd__decap_3 PHY_1649 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_1650 ();
 sky130_fd_sc_hd__decap_3 PHY_1651 ();
 sky130_fd_sc_hd__decap_3 PHY_1652 ();
 sky130_fd_sc_hd__decap_3 PHY_1653 ();
 sky130_fd_sc_hd__decap_3 PHY_1654 ();
 sky130_fd_sc_hd__decap_3 PHY_1655 ();
 sky130_fd_sc_hd__decap_3 PHY_1656 ();
 sky130_fd_sc_hd__decap_3 PHY_1657 ();
 sky130_fd_sc_hd__decap_3 PHY_1658 ();
 sky130_fd_sc_hd__decap_3 PHY_1659 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_1660 ();
 sky130_fd_sc_hd__decap_3 PHY_1661 ();
 sky130_fd_sc_hd__decap_3 PHY_1662 ();
 sky130_fd_sc_hd__decap_3 PHY_1663 ();
 sky130_fd_sc_hd__decap_3 PHY_1664 ();
 sky130_fd_sc_hd__decap_3 PHY_1665 ();
 sky130_fd_sc_hd__decap_3 PHY_1666 ();
 sky130_fd_sc_hd__decap_3 PHY_1667 ();
 sky130_fd_sc_hd__decap_3 PHY_1668 ();
 sky130_fd_sc_hd__decap_3 PHY_1669 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_1670 ();
 sky130_fd_sc_hd__decap_3 PHY_1671 ();
 sky130_fd_sc_hd__decap_3 PHY_1672 ();
 sky130_fd_sc_hd__decap_3 PHY_1673 ();
 sky130_fd_sc_hd__decap_3 PHY_1674 ();
 sky130_fd_sc_hd__decap_3 PHY_1675 ();
 sky130_fd_sc_hd__decap_3 PHY_1676 ();
 sky130_fd_sc_hd__decap_3 PHY_1677 ();
 sky130_fd_sc_hd__decap_3 PHY_1678 ();
 sky130_fd_sc_hd__decap_3 PHY_1679 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_1680 ();
 sky130_fd_sc_hd__decap_3 PHY_1681 ();
 sky130_fd_sc_hd__decap_3 PHY_1682 ();
 sky130_fd_sc_hd__decap_3 PHY_1683 ();
 sky130_fd_sc_hd__decap_3 PHY_1684 ();
 sky130_fd_sc_hd__decap_3 PHY_1685 ();
 sky130_fd_sc_hd__decap_3 PHY_1686 ();
 sky130_fd_sc_hd__decap_3 PHY_1687 ();
 sky130_fd_sc_hd__decap_3 PHY_1688 ();
 sky130_fd_sc_hd__decap_3 PHY_1689 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_1690 ();
 sky130_fd_sc_hd__decap_3 PHY_1691 ();
 sky130_fd_sc_hd__decap_3 PHY_1692 ();
 sky130_fd_sc_hd__decap_3 PHY_1693 ();
 sky130_fd_sc_hd__decap_3 PHY_1694 ();
 sky130_fd_sc_hd__decap_3 PHY_1695 ();
 sky130_fd_sc_hd__decap_3 PHY_1696 ();
 sky130_fd_sc_hd__decap_3 PHY_1697 ();
 sky130_fd_sc_hd__decap_3 PHY_1698 ();
 sky130_fd_sc_hd__decap_3 PHY_1699 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_1700 ();
 sky130_fd_sc_hd__decap_3 PHY_1701 ();
 sky130_fd_sc_hd__decap_3 PHY_1702 ();
 sky130_fd_sc_hd__decap_3 PHY_1703 ();
 sky130_fd_sc_hd__decap_3 PHY_1704 ();
 sky130_fd_sc_hd__decap_3 PHY_1705 ();
 sky130_fd_sc_hd__decap_3 PHY_1706 ();
 sky130_fd_sc_hd__decap_3 PHY_1707 ();
 sky130_fd_sc_hd__decap_3 PHY_1708 ();
 sky130_fd_sc_hd__decap_3 PHY_1709 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_1710 ();
 sky130_fd_sc_hd__decap_3 PHY_1711 ();
 sky130_fd_sc_hd__decap_3 PHY_1712 ();
 sky130_fd_sc_hd__decap_3 PHY_1713 ();
 sky130_fd_sc_hd__decap_3 PHY_1714 ();
 sky130_fd_sc_hd__decap_3 PHY_1715 ();
 sky130_fd_sc_hd__decap_3 PHY_1716 ();
 sky130_fd_sc_hd__decap_3 PHY_1717 ();
 sky130_fd_sc_hd__decap_3 PHY_1718 ();
 sky130_fd_sc_hd__decap_3 PHY_1719 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_1720 ();
 sky130_fd_sc_hd__decap_3 PHY_1721 ();
 sky130_fd_sc_hd__decap_3 PHY_1722 ();
 sky130_fd_sc_hd__decap_3 PHY_1723 ();
 sky130_fd_sc_hd__decap_3 PHY_1724 ();
 sky130_fd_sc_hd__decap_3 PHY_1725 ();
 sky130_fd_sc_hd__decap_3 PHY_1726 ();
 sky130_fd_sc_hd__decap_3 PHY_1727 ();
 sky130_fd_sc_hd__decap_3 PHY_1728 ();
 sky130_fd_sc_hd__decap_3 PHY_1729 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_1730 ();
 sky130_fd_sc_hd__decap_3 PHY_1731 ();
 sky130_fd_sc_hd__decap_3 PHY_1732 ();
 sky130_fd_sc_hd__decap_3 PHY_1733 ();
 sky130_fd_sc_hd__decap_3 PHY_1734 ();
 sky130_fd_sc_hd__decap_3 PHY_1735 ();
 sky130_fd_sc_hd__decap_3 PHY_1736 ();
 sky130_fd_sc_hd__decap_3 PHY_1737 ();
 sky130_fd_sc_hd__decap_3 PHY_1738 ();
 sky130_fd_sc_hd__decap_3 PHY_1739 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_1740 ();
 sky130_fd_sc_hd__decap_3 PHY_1741 ();
 sky130_fd_sc_hd__decap_3 PHY_1742 ();
 sky130_fd_sc_hd__decap_3 PHY_1743 ();
 sky130_fd_sc_hd__decap_3 PHY_1744 ();
 sky130_fd_sc_hd__decap_3 PHY_1745 ();
 sky130_fd_sc_hd__decap_3 PHY_1746 ();
 sky130_fd_sc_hd__decap_3 PHY_1747 ();
 sky130_fd_sc_hd__decap_3 PHY_1748 ();
 sky130_fd_sc_hd__decap_3 PHY_1749 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_1750 ();
 sky130_fd_sc_hd__decap_3 PHY_1751 ();
 sky130_fd_sc_hd__decap_3 PHY_1752 ();
 sky130_fd_sc_hd__decap_3 PHY_1753 ();
 sky130_fd_sc_hd__decap_3 PHY_1754 ();
 sky130_fd_sc_hd__decap_3 PHY_1755 ();
 sky130_fd_sc_hd__decap_3 PHY_1756 ();
 sky130_fd_sc_hd__decap_3 PHY_1757 ();
 sky130_fd_sc_hd__decap_3 PHY_1758 ();
 sky130_fd_sc_hd__decap_3 PHY_1759 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_1760 ();
 sky130_fd_sc_hd__decap_3 PHY_1761 ();
 sky130_fd_sc_hd__decap_3 PHY_1762 ();
 sky130_fd_sc_hd__decap_3 PHY_1763 ();
 sky130_fd_sc_hd__decap_3 PHY_1764 ();
 sky130_fd_sc_hd__decap_3 PHY_1765 ();
 sky130_fd_sc_hd__decap_3 PHY_1766 ();
 sky130_fd_sc_hd__decap_3 PHY_1767 ();
 sky130_fd_sc_hd__decap_3 PHY_1768 ();
 sky130_fd_sc_hd__decap_3 PHY_1769 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_1770 ();
 sky130_fd_sc_hd__decap_3 PHY_1771 ();
 sky130_fd_sc_hd__decap_3 PHY_1772 ();
 sky130_fd_sc_hd__decap_3 PHY_1773 ();
 sky130_fd_sc_hd__decap_3 PHY_1774 ();
 sky130_fd_sc_hd__decap_3 PHY_1775 ();
 sky130_fd_sc_hd__decap_3 PHY_1776 ();
 sky130_fd_sc_hd__decap_3 PHY_1777 ();
 sky130_fd_sc_hd__decap_3 PHY_1778 ();
 sky130_fd_sc_hd__decap_3 PHY_1779 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_1780 ();
 sky130_fd_sc_hd__decap_3 PHY_1781 ();
 sky130_fd_sc_hd__decap_3 PHY_1782 ();
 sky130_fd_sc_hd__decap_3 PHY_1783 ();
 sky130_fd_sc_hd__decap_3 PHY_1784 ();
 sky130_fd_sc_hd__decap_3 PHY_1785 ();
 sky130_fd_sc_hd__decap_3 PHY_1786 ();
 sky130_fd_sc_hd__decap_3 PHY_1787 ();
 sky130_fd_sc_hd__decap_3 PHY_1788 ();
 sky130_fd_sc_hd__decap_3 PHY_1789 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_1790 ();
 sky130_fd_sc_hd__decap_3 PHY_1791 ();
 sky130_fd_sc_hd__decap_3 PHY_1792 ();
 sky130_fd_sc_hd__decap_3 PHY_1793 ();
 sky130_fd_sc_hd__decap_3 PHY_1794 ();
 sky130_fd_sc_hd__decap_3 PHY_1795 ();
 sky130_fd_sc_hd__decap_3 PHY_1796 ();
 sky130_fd_sc_hd__decap_3 PHY_1797 ();
 sky130_fd_sc_hd__decap_3 PHY_1798 ();
 sky130_fd_sc_hd__decap_3 PHY_1799 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_1800 ();
 sky130_fd_sc_hd__decap_3 PHY_1801 ();
 sky130_fd_sc_hd__decap_3 PHY_1802 ();
 sky130_fd_sc_hd__decap_3 PHY_1803 ();
 sky130_fd_sc_hd__decap_3 PHY_1804 ();
 sky130_fd_sc_hd__decap_3 PHY_1805 ();
 sky130_fd_sc_hd__decap_3 PHY_1806 ();
 sky130_fd_sc_hd__decap_3 PHY_1807 ();
 sky130_fd_sc_hd__decap_3 PHY_1808 ();
 sky130_fd_sc_hd__decap_3 PHY_1809 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_1810 ();
 sky130_fd_sc_hd__decap_3 PHY_1811 ();
 sky130_fd_sc_hd__decap_3 PHY_1812 ();
 sky130_fd_sc_hd__decap_3 PHY_1813 ();
 sky130_fd_sc_hd__decap_3 PHY_1814 ();
 sky130_fd_sc_hd__decap_3 PHY_1815 ();
 sky130_fd_sc_hd__decap_3 PHY_1816 ();
 sky130_fd_sc_hd__decap_3 PHY_1817 ();
 sky130_fd_sc_hd__decap_3 PHY_1818 ();
 sky130_fd_sc_hd__decap_3 PHY_1819 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_1820 ();
 sky130_fd_sc_hd__decap_3 PHY_1821 ();
 sky130_fd_sc_hd__decap_3 PHY_1822 ();
 sky130_fd_sc_hd__decap_3 PHY_1823 ();
 sky130_fd_sc_hd__decap_3 PHY_1824 ();
 sky130_fd_sc_hd__decap_3 PHY_1825 ();
 sky130_fd_sc_hd__decap_3 PHY_1826 ();
 sky130_fd_sc_hd__decap_3 PHY_1827 ();
 sky130_fd_sc_hd__decap_3 PHY_1828 ();
 sky130_fd_sc_hd__decap_3 PHY_1829 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_1830 ();
 sky130_fd_sc_hd__decap_3 PHY_1831 ();
 sky130_fd_sc_hd__decap_3 PHY_1832 ();
 sky130_fd_sc_hd__decap_3 PHY_1833 ();
 sky130_fd_sc_hd__decap_3 PHY_1834 ();
 sky130_fd_sc_hd__decap_3 PHY_1835 ();
 sky130_fd_sc_hd__decap_3 PHY_1836 ();
 sky130_fd_sc_hd__decap_3 PHY_1837 ();
 sky130_fd_sc_hd__decap_3 PHY_1838 ();
 sky130_fd_sc_hd__decap_3 PHY_1839 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_1840 ();
 sky130_fd_sc_hd__decap_3 PHY_1841 ();
 sky130_fd_sc_hd__decap_3 PHY_1842 ();
 sky130_fd_sc_hd__decap_3 PHY_1843 ();
 sky130_fd_sc_hd__decap_3 PHY_1844 ();
 sky130_fd_sc_hd__decap_3 PHY_1845 ();
 sky130_fd_sc_hd__decap_3 PHY_1846 ();
 sky130_fd_sc_hd__decap_3 PHY_1847 ();
 sky130_fd_sc_hd__decap_3 PHY_1848 ();
 sky130_fd_sc_hd__decap_3 PHY_1849 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_1850 ();
 sky130_fd_sc_hd__decap_3 PHY_1851 ();
 sky130_fd_sc_hd__decap_3 PHY_1852 ();
 sky130_fd_sc_hd__decap_3 PHY_1853 ();
 sky130_fd_sc_hd__decap_3 PHY_1854 ();
 sky130_fd_sc_hd__decap_3 PHY_1855 ();
 sky130_fd_sc_hd__decap_3 PHY_1856 ();
 sky130_fd_sc_hd__decap_3 PHY_1857 ();
 sky130_fd_sc_hd__decap_3 PHY_1858 ();
 sky130_fd_sc_hd__decap_3 PHY_1859 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_1860 ();
 sky130_fd_sc_hd__decap_3 PHY_1861 ();
 sky130_fd_sc_hd__decap_3 PHY_1862 ();
 sky130_fd_sc_hd__decap_3 PHY_1863 ();
 sky130_fd_sc_hd__decap_3 PHY_1864 ();
 sky130_fd_sc_hd__decap_3 PHY_1865 ();
 sky130_fd_sc_hd__decap_3 PHY_1866 ();
 sky130_fd_sc_hd__decap_3 PHY_1867 ();
 sky130_fd_sc_hd__decap_3 PHY_1868 ();
 sky130_fd_sc_hd__decap_3 PHY_1869 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_1870 ();
 sky130_fd_sc_hd__decap_3 PHY_1871 ();
 sky130_fd_sc_hd__decap_3 PHY_1872 ();
 sky130_fd_sc_hd__decap_3 PHY_1873 ();
 sky130_fd_sc_hd__decap_3 PHY_1874 ();
 sky130_fd_sc_hd__decap_3 PHY_1875 ();
 sky130_fd_sc_hd__decap_3 PHY_1876 ();
 sky130_fd_sc_hd__decap_3 PHY_1877 ();
 sky130_fd_sc_hd__decap_3 PHY_1878 ();
 sky130_fd_sc_hd__decap_3 PHY_1879 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_1880 ();
 sky130_fd_sc_hd__decap_3 PHY_1881 ();
 sky130_fd_sc_hd__decap_3 PHY_1882 ();
 sky130_fd_sc_hd__decap_3 PHY_1883 ();
 sky130_fd_sc_hd__decap_3 PHY_1884 ();
 sky130_fd_sc_hd__decap_3 PHY_1885 ();
 sky130_fd_sc_hd__decap_3 PHY_1886 ();
 sky130_fd_sc_hd__decap_3 PHY_1887 ();
 sky130_fd_sc_hd__decap_3 PHY_1888 ();
 sky130_fd_sc_hd__decap_3 PHY_1889 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_1890 ();
 sky130_fd_sc_hd__decap_3 PHY_1891 ();
 sky130_fd_sc_hd__decap_3 PHY_1892 ();
 sky130_fd_sc_hd__decap_3 PHY_1893 ();
 sky130_fd_sc_hd__decap_3 PHY_1894 ();
 sky130_fd_sc_hd__decap_3 PHY_1895 ();
 sky130_fd_sc_hd__decap_3 PHY_1896 ();
 sky130_fd_sc_hd__decap_3 PHY_1897 ();
 sky130_fd_sc_hd__decap_3 PHY_1898 ();
 sky130_fd_sc_hd__decap_3 PHY_1899 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_1900 ();
 sky130_fd_sc_hd__decap_3 PHY_1901 ();
 sky130_fd_sc_hd__decap_3 PHY_1902 ();
 sky130_fd_sc_hd__decap_3 PHY_1903 ();
 sky130_fd_sc_hd__decap_3 PHY_1904 ();
 sky130_fd_sc_hd__decap_3 PHY_1905 ();
 sky130_fd_sc_hd__decap_3 PHY_1906 ();
 sky130_fd_sc_hd__decap_3 PHY_1907 ();
 sky130_fd_sc_hd__decap_3 PHY_1908 ();
 sky130_fd_sc_hd__decap_3 PHY_1909 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_1910 ();
 sky130_fd_sc_hd__decap_3 PHY_1911 ();
 sky130_fd_sc_hd__decap_3 PHY_1912 ();
 sky130_fd_sc_hd__decap_3 PHY_1913 ();
 sky130_fd_sc_hd__decap_3 PHY_1914 ();
 sky130_fd_sc_hd__decap_3 PHY_1915 ();
 sky130_fd_sc_hd__decap_3 PHY_1916 ();
 sky130_fd_sc_hd__decap_3 PHY_1917 ();
 sky130_fd_sc_hd__decap_3 PHY_1918 ();
 sky130_fd_sc_hd__decap_3 PHY_1919 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_1920 ();
 sky130_fd_sc_hd__decap_3 PHY_1921 ();
 sky130_fd_sc_hd__decap_3 PHY_1922 ();
 sky130_fd_sc_hd__decap_3 PHY_1923 ();
 sky130_fd_sc_hd__decap_3 PHY_1924 ();
 sky130_fd_sc_hd__decap_3 PHY_1925 ();
 sky130_fd_sc_hd__decap_3 PHY_1926 ();
 sky130_fd_sc_hd__decap_3 PHY_1927 ();
 sky130_fd_sc_hd__decap_3 PHY_1928 ();
 sky130_fd_sc_hd__decap_3 PHY_1929 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_1930 ();
 sky130_fd_sc_hd__decap_3 PHY_1931 ();
 sky130_fd_sc_hd__decap_3 PHY_1932 ();
 sky130_fd_sc_hd__decap_3 PHY_1933 ();
 sky130_fd_sc_hd__decap_3 PHY_1934 ();
 sky130_fd_sc_hd__decap_3 PHY_1935 ();
 sky130_fd_sc_hd__decap_3 PHY_1936 ();
 sky130_fd_sc_hd__decap_3 PHY_1937 ();
 sky130_fd_sc_hd__decap_3 PHY_1938 ();
 sky130_fd_sc_hd__decap_3 PHY_1939 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_1940 ();
 sky130_fd_sc_hd__decap_3 PHY_1941 ();
 sky130_fd_sc_hd__decap_3 PHY_1942 ();
 sky130_fd_sc_hd__decap_3 PHY_1943 ();
 sky130_fd_sc_hd__decap_3 PHY_1944 ();
 sky130_fd_sc_hd__decap_3 PHY_1945 ();
 sky130_fd_sc_hd__decap_3 PHY_1946 ();
 sky130_fd_sc_hd__decap_3 PHY_1947 ();
 sky130_fd_sc_hd__decap_3 PHY_1948 ();
 sky130_fd_sc_hd__decap_3 PHY_1949 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_1950 ();
 sky130_fd_sc_hd__decap_3 PHY_1951 ();
 sky130_fd_sc_hd__decap_3 PHY_1952 ();
 sky130_fd_sc_hd__decap_3 PHY_1953 ();
 sky130_fd_sc_hd__decap_3 PHY_1954 ();
 sky130_fd_sc_hd__decap_3 PHY_1955 ();
 sky130_fd_sc_hd__decap_3 PHY_1956 ();
 sky130_fd_sc_hd__decap_3 PHY_1957 ();
 sky130_fd_sc_hd__decap_3 PHY_1958 ();
 sky130_fd_sc_hd__decap_3 PHY_1959 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_1960 ();
 sky130_fd_sc_hd__decap_3 PHY_1961 ();
 sky130_fd_sc_hd__decap_3 PHY_1962 ();
 sky130_fd_sc_hd__decap_3 PHY_1963 ();
 sky130_fd_sc_hd__decap_3 PHY_1964 ();
 sky130_fd_sc_hd__decap_3 PHY_1965 ();
 sky130_fd_sc_hd__decap_3 PHY_1966 ();
 sky130_fd_sc_hd__decap_3 PHY_1967 ();
 sky130_fd_sc_hd__decap_3 PHY_1968 ();
 sky130_fd_sc_hd__decap_3 PHY_1969 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_1970 ();
 sky130_fd_sc_hd__decap_3 PHY_1971 ();
 sky130_fd_sc_hd__decap_3 PHY_1972 ();
 sky130_fd_sc_hd__decap_3 PHY_1973 ();
 sky130_fd_sc_hd__decap_3 PHY_1974 ();
 sky130_fd_sc_hd__decap_3 PHY_1975 ();
 sky130_fd_sc_hd__decap_3 PHY_1976 ();
 sky130_fd_sc_hd__decap_3 PHY_1977 ();
 sky130_fd_sc_hd__decap_3 PHY_1978 ();
 sky130_fd_sc_hd__decap_3 PHY_1979 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_1980 ();
 sky130_fd_sc_hd__decap_3 PHY_1981 ();
 sky130_fd_sc_hd__decap_3 PHY_1982 ();
 sky130_fd_sc_hd__decap_3 PHY_1983 ();
 sky130_fd_sc_hd__decap_3 PHY_1984 ();
 sky130_fd_sc_hd__decap_3 PHY_1985 ();
 sky130_fd_sc_hd__decap_3 PHY_1986 ();
 sky130_fd_sc_hd__decap_3 PHY_1987 ();
 sky130_fd_sc_hd__decap_3 PHY_1988 ();
 sky130_fd_sc_hd__decap_3 PHY_1989 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_1990 ();
 sky130_fd_sc_hd__decap_3 PHY_1991 ();
 sky130_fd_sc_hd__decap_3 PHY_1992 ();
 sky130_fd_sc_hd__decap_3 PHY_1993 ();
 sky130_fd_sc_hd__decap_3 PHY_1994 ();
 sky130_fd_sc_hd__decap_3 PHY_1995 ();
 sky130_fd_sc_hd__decap_3 PHY_1996 ();
 sky130_fd_sc_hd__decap_3 PHY_1997 ();
 sky130_fd_sc_hd__decap_3 PHY_1998 ();
 sky130_fd_sc_hd__decap_3 PHY_1999 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_2000 ();
 sky130_fd_sc_hd__decap_3 PHY_2001 ();
 sky130_fd_sc_hd__decap_3 PHY_2002 ();
 sky130_fd_sc_hd__decap_3 PHY_2003 ();
 sky130_fd_sc_hd__decap_3 PHY_2004 ();
 sky130_fd_sc_hd__decap_3 PHY_2005 ();
 sky130_fd_sc_hd__decap_3 PHY_2006 ();
 sky130_fd_sc_hd__decap_3 PHY_2007 ();
 sky130_fd_sc_hd__decap_3 PHY_2008 ();
 sky130_fd_sc_hd__decap_3 PHY_2009 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_2010 ();
 sky130_fd_sc_hd__decap_3 PHY_2011 ();
 sky130_fd_sc_hd__decap_3 PHY_2012 ();
 sky130_fd_sc_hd__decap_3 PHY_2013 ();
 sky130_fd_sc_hd__decap_3 PHY_2014 ();
 sky130_fd_sc_hd__decap_3 PHY_2015 ();
 sky130_fd_sc_hd__decap_3 PHY_2016 ();
 sky130_fd_sc_hd__decap_3 PHY_2017 ();
 sky130_fd_sc_hd__decap_3 PHY_2018 ();
 sky130_fd_sc_hd__decap_3 PHY_2019 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_2020 ();
 sky130_fd_sc_hd__decap_3 PHY_2021 ();
 sky130_fd_sc_hd__decap_3 PHY_2022 ();
 sky130_fd_sc_hd__decap_3 PHY_2023 ();
 sky130_fd_sc_hd__decap_3 PHY_2024 ();
 sky130_fd_sc_hd__decap_3 PHY_2025 ();
 sky130_fd_sc_hd__decap_3 PHY_2026 ();
 sky130_fd_sc_hd__decap_3 PHY_2027 ();
 sky130_fd_sc_hd__decap_3 PHY_2028 ();
 sky130_fd_sc_hd__decap_3 PHY_2029 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_2030 ();
 sky130_fd_sc_hd__decap_3 PHY_2031 ();
 sky130_fd_sc_hd__decap_3 PHY_2032 ();
 sky130_fd_sc_hd__decap_3 PHY_2033 ();
 sky130_fd_sc_hd__decap_3 PHY_2034 ();
 sky130_fd_sc_hd__decap_3 PHY_2035 ();
 sky130_fd_sc_hd__decap_3 PHY_2036 ();
 sky130_fd_sc_hd__decap_3 PHY_2037 ();
 sky130_fd_sc_hd__decap_3 PHY_2038 ();
 sky130_fd_sc_hd__decap_3 PHY_2039 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_2040 ();
 sky130_fd_sc_hd__decap_3 PHY_2041 ();
 sky130_fd_sc_hd__decap_3 PHY_2042 ();
 sky130_fd_sc_hd__decap_3 PHY_2043 ();
 sky130_fd_sc_hd__decap_3 PHY_2044 ();
 sky130_fd_sc_hd__decap_3 PHY_2045 ();
 sky130_fd_sc_hd__decap_3 PHY_2046 ();
 sky130_fd_sc_hd__decap_3 PHY_2047 ();
 sky130_fd_sc_hd__decap_3 PHY_2048 ();
 sky130_fd_sc_hd__decap_3 PHY_2049 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_2050 ();
 sky130_fd_sc_hd__decap_3 PHY_2051 ();
 sky130_fd_sc_hd__decap_3 PHY_2052 ();
 sky130_fd_sc_hd__decap_3 PHY_2053 ();
 sky130_fd_sc_hd__decap_3 PHY_2054 ();
 sky130_fd_sc_hd__decap_3 PHY_2055 ();
 sky130_fd_sc_hd__decap_3 PHY_2056 ();
 sky130_fd_sc_hd__decap_3 PHY_2057 ();
 sky130_fd_sc_hd__decap_3 PHY_2058 ();
 sky130_fd_sc_hd__decap_3 PHY_2059 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_2060 ();
 sky130_fd_sc_hd__decap_3 PHY_2061 ();
 sky130_fd_sc_hd__decap_3 PHY_2062 ();
 sky130_fd_sc_hd__decap_3 PHY_2063 ();
 sky130_fd_sc_hd__decap_3 PHY_2064 ();
 sky130_fd_sc_hd__decap_3 PHY_2065 ();
 sky130_fd_sc_hd__decap_3 PHY_2066 ();
 sky130_fd_sc_hd__decap_3 PHY_2067 ();
 sky130_fd_sc_hd__decap_3 PHY_2068 ();
 sky130_fd_sc_hd__decap_3 PHY_2069 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_2070 ();
 sky130_fd_sc_hd__decap_3 PHY_2071 ();
 sky130_fd_sc_hd__decap_3 PHY_2072 ();
 sky130_fd_sc_hd__decap_3 PHY_2073 ();
 sky130_fd_sc_hd__decap_3 PHY_2074 ();
 sky130_fd_sc_hd__decap_3 PHY_2075 ();
 sky130_fd_sc_hd__decap_3 PHY_2076 ();
 sky130_fd_sc_hd__decap_3 PHY_2077 ();
 sky130_fd_sc_hd__decap_3 PHY_2078 ();
 sky130_fd_sc_hd__decap_3 PHY_2079 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_2080 ();
 sky130_fd_sc_hd__decap_3 PHY_2081 ();
 sky130_fd_sc_hd__decap_3 PHY_2082 ();
 sky130_fd_sc_hd__decap_3 PHY_2083 ();
 sky130_fd_sc_hd__decap_3 PHY_2084 ();
 sky130_fd_sc_hd__decap_3 PHY_2085 ();
 sky130_fd_sc_hd__decap_3 PHY_2086 ();
 sky130_fd_sc_hd__decap_3 PHY_2087 ();
 sky130_fd_sc_hd__decap_3 PHY_2088 ();
 sky130_fd_sc_hd__decap_3 PHY_2089 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_2090 ();
 sky130_fd_sc_hd__decap_3 PHY_2091 ();
 sky130_fd_sc_hd__decap_3 PHY_2092 ();
 sky130_fd_sc_hd__decap_3 PHY_2093 ();
 sky130_fd_sc_hd__decap_3 PHY_2094 ();
 sky130_fd_sc_hd__decap_3 PHY_2095 ();
 sky130_fd_sc_hd__decap_3 PHY_2096 ();
 sky130_fd_sc_hd__decap_3 PHY_2097 ();
 sky130_fd_sc_hd__decap_3 PHY_2098 ();
 sky130_fd_sc_hd__decap_3 PHY_2099 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_2100 ();
 sky130_fd_sc_hd__decap_3 PHY_2101 ();
 sky130_fd_sc_hd__decap_3 PHY_2102 ();
 sky130_fd_sc_hd__decap_3 PHY_2103 ();
 sky130_fd_sc_hd__decap_3 PHY_2104 ();
 sky130_fd_sc_hd__decap_3 PHY_2105 ();
 sky130_fd_sc_hd__decap_3 PHY_2106 ();
 sky130_fd_sc_hd__decap_3 PHY_2107 ();
 sky130_fd_sc_hd__decap_3 PHY_2108 ();
 sky130_fd_sc_hd__decap_3 PHY_2109 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_2110 ();
 sky130_fd_sc_hd__decap_3 PHY_2111 ();
 sky130_fd_sc_hd__decap_3 PHY_2112 ();
 sky130_fd_sc_hd__decap_3 PHY_2113 ();
 sky130_fd_sc_hd__decap_3 PHY_2114 ();
 sky130_fd_sc_hd__decap_3 PHY_2115 ();
 sky130_fd_sc_hd__decap_3 PHY_2116 ();
 sky130_fd_sc_hd__decap_3 PHY_2117 ();
 sky130_fd_sc_hd__decap_3 PHY_2118 ();
 sky130_fd_sc_hd__decap_3 PHY_2119 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_2120 ();
 sky130_fd_sc_hd__decap_3 PHY_2121 ();
 sky130_fd_sc_hd__decap_3 PHY_2122 ();
 sky130_fd_sc_hd__decap_3 PHY_2123 ();
 sky130_fd_sc_hd__decap_3 PHY_2124 ();
 sky130_fd_sc_hd__decap_3 PHY_2125 ();
 sky130_fd_sc_hd__decap_3 PHY_2126 ();
 sky130_fd_sc_hd__decap_3 PHY_2127 ();
 sky130_fd_sc_hd__decap_3 PHY_2128 ();
 sky130_fd_sc_hd__decap_3 PHY_2129 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_2130 ();
 sky130_fd_sc_hd__decap_3 PHY_2131 ();
 sky130_fd_sc_hd__decap_3 PHY_2132 ();
 sky130_fd_sc_hd__decap_3 PHY_2133 ();
 sky130_fd_sc_hd__decap_3 PHY_2134 ();
 sky130_fd_sc_hd__decap_3 PHY_2135 ();
 sky130_fd_sc_hd__decap_3 PHY_2136 ();
 sky130_fd_sc_hd__decap_3 PHY_2137 ();
 sky130_fd_sc_hd__decap_3 PHY_2138 ();
 sky130_fd_sc_hd__decap_3 PHY_2139 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_2140 ();
 sky130_fd_sc_hd__decap_3 PHY_2141 ();
 sky130_fd_sc_hd__decap_3 PHY_2142 ();
 sky130_fd_sc_hd__decap_3 PHY_2143 ();
 sky130_fd_sc_hd__decap_3 PHY_2144 ();
 sky130_fd_sc_hd__decap_3 PHY_2145 ();
 sky130_fd_sc_hd__decap_3 PHY_2146 ();
 sky130_fd_sc_hd__decap_3 PHY_2147 ();
 sky130_fd_sc_hd__decap_3 PHY_2148 ();
 sky130_fd_sc_hd__decap_3 PHY_2149 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_2150 ();
 sky130_fd_sc_hd__decap_3 PHY_2151 ();
 sky130_fd_sc_hd__decap_3 PHY_2152 ();
 sky130_fd_sc_hd__decap_3 PHY_2153 ();
 sky130_fd_sc_hd__decap_3 PHY_2154 ();
 sky130_fd_sc_hd__decap_3 PHY_2155 ();
 sky130_fd_sc_hd__decap_3 PHY_2156 ();
 sky130_fd_sc_hd__decap_3 PHY_2157 ();
 sky130_fd_sc_hd__decap_3 PHY_2158 ();
 sky130_fd_sc_hd__decap_3 PHY_2159 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_2160 ();
 sky130_fd_sc_hd__decap_3 PHY_2161 ();
 sky130_fd_sc_hd__decap_3 PHY_2162 ();
 sky130_fd_sc_hd__decap_3 PHY_2163 ();
 sky130_fd_sc_hd__decap_3 PHY_2164 ();
 sky130_fd_sc_hd__decap_3 PHY_2165 ();
 sky130_fd_sc_hd__decap_3 PHY_2166 ();
 sky130_fd_sc_hd__decap_3 PHY_2167 ();
 sky130_fd_sc_hd__decap_3 PHY_2168 ();
 sky130_fd_sc_hd__decap_3 PHY_2169 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_2170 ();
 sky130_fd_sc_hd__decap_3 PHY_2171 ();
 sky130_fd_sc_hd__decap_3 PHY_2172 ();
 sky130_fd_sc_hd__decap_3 PHY_2173 ();
 sky130_fd_sc_hd__decap_3 PHY_2174 ();
 sky130_fd_sc_hd__decap_3 PHY_2175 ();
 sky130_fd_sc_hd__decap_3 PHY_2176 ();
 sky130_fd_sc_hd__decap_3 PHY_2177 ();
 sky130_fd_sc_hd__decap_3 PHY_2178 ();
 sky130_fd_sc_hd__decap_3 PHY_2179 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_2180 ();
 sky130_fd_sc_hd__decap_3 PHY_2181 ();
 sky130_fd_sc_hd__decap_3 PHY_2182 ();
 sky130_fd_sc_hd__decap_3 PHY_2183 ();
 sky130_fd_sc_hd__decap_3 PHY_2184 ();
 sky130_fd_sc_hd__decap_3 PHY_2185 ();
 sky130_fd_sc_hd__decap_3 PHY_2186 ();
 sky130_fd_sc_hd__decap_3 PHY_2187 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_880 ();
 sky130_fd_sc_hd__decap_3 PHY_881 ();
 sky130_fd_sc_hd__decap_3 PHY_882 ();
 sky130_fd_sc_hd__decap_3 PHY_883 ();
 sky130_fd_sc_hd__decap_3 PHY_884 ();
 sky130_fd_sc_hd__decap_3 PHY_885 ();
 sky130_fd_sc_hd__decap_3 PHY_886 ();
 sky130_fd_sc_hd__decap_3 PHY_887 ();
 sky130_fd_sc_hd__decap_3 PHY_888 ();
 sky130_fd_sc_hd__decap_3 PHY_889 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_890 ();
 sky130_fd_sc_hd__decap_3 PHY_891 ();
 sky130_fd_sc_hd__decap_3 PHY_892 ();
 sky130_fd_sc_hd__decap_3 PHY_893 ();
 sky130_fd_sc_hd__decap_3 PHY_894 ();
 sky130_fd_sc_hd__decap_3 PHY_895 ();
 sky130_fd_sc_hd__decap_3 PHY_896 ();
 sky130_fd_sc_hd__decap_3 PHY_897 ();
 sky130_fd_sc_hd__decap_3 PHY_898 ();
 sky130_fd_sc_hd__decap_3 PHY_899 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_900 ();
 sky130_fd_sc_hd__decap_3 PHY_901 ();
 sky130_fd_sc_hd__decap_3 PHY_902 ();
 sky130_fd_sc_hd__decap_3 PHY_903 ();
 sky130_fd_sc_hd__decap_3 PHY_904 ();
 sky130_fd_sc_hd__decap_3 PHY_905 ();
 sky130_fd_sc_hd__decap_3 PHY_906 ();
 sky130_fd_sc_hd__decap_3 PHY_907 ();
 sky130_fd_sc_hd__decap_3 PHY_908 ();
 sky130_fd_sc_hd__decap_3 PHY_909 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_910 ();
 sky130_fd_sc_hd__decap_3 PHY_911 ();
 sky130_fd_sc_hd__decap_3 PHY_912 ();
 sky130_fd_sc_hd__decap_3 PHY_913 ();
 sky130_fd_sc_hd__decap_3 PHY_914 ();
 sky130_fd_sc_hd__decap_3 PHY_915 ();
 sky130_fd_sc_hd__decap_3 PHY_916 ();
 sky130_fd_sc_hd__decap_3 PHY_917 ();
 sky130_fd_sc_hd__decap_3 PHY_918 ();
 sky130_fd_sc_hd__decap_3 PHY_919 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_920 ();
 sky130_fd_sc_hd__decap_3 PHY_921 ();
 sky130_fd_sc_hd__decap_3 PHY_922 ();
 sky130_fd_sc_hd__decap_3 PHY_923 ();
 sky130_fd_sc_hd__decap_3 PHY_924 ();
 sky130_fd_sc_hd__decap_3 PHY_925 ();
 sky130_fd_sc_hd__decap_3 PHY_926 ();
 sky130_fd_sc_hd__decap_3 PHY_927 ();
 sky130_fd_sc_hd__decap_3 PHY_928 ();
 sky130_fd_sc_hd__decap_3 PHY_929 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_930 ();
 sky130_fd_sc_hd__decap_3 PHY_931 ();
 sky130_fd_sc_hd__decap_3 PHY_932 ();
 sky130_fd_sc_hd__decap_3 PHY_933 ();
 sky130_fd_sc_hd__decap_3 PHY_934 ();
 sky130_fd_sc_hd__decap_3 PHY_935 ();
 sky130_fd_sc_hd__decap_3 PHY_936 ();
 sky130_fd_sc_hd__decap_3 PHY_937 ();
 sky130_fd_sc_hd__decap_3 PHY_938 ();
 sky130_fd_sc_hd__decap_3 PHY_939 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_940 ();
 sky130_fd_sc_hd__decap_3 PHY_941 ();
 sky130_fd_sc_hd__decap_3 PHY_942 ();
 sky130_fd_sc_hd__decap_3 PHY_943 ();
 sky130_fd_sc_hd__decap_3 PHY_944 ();
 sky130_fd_sc_hd__decap_3 PHY_945 ();
 sky130_fd_sc_hd__decap_3 PHY_946 ();
 sky130_fd_sc_hd__decap_3 PHY_947 ();
 sky130_fd_sc_hd__decap_3 PHY_948 ();
 sky130_fd_sc_hd__decap_3 PHY_949 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_950 ();
 sky130_fd_sc_hd__decap_3 PHY_951 ();
 sky130_fd_sc_hd__decap_3 PHY_952 ();
 sky130_fd_sc_hd__decap_3 PHY_953 ();
 sky130_fd_sc_hd__decap_3 PHY_954 ();
 sky130_fd_sc_hd__decap_3 PHY_955 ();
 sky130_fd_sc_hd__decap_3 PHY_956 ();
 sky130_fd_sc_hd__decap_3 PHY_957 ();
 sky130_fd_sc_hd__decap_3 PHY_958 ();
 sky130_fd_sc_hd__decap_3 PHY_959 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_960 ();
 sky130_fd_sc_hd__decap_3 PHY_961 ();
 sky130_fd_sc_hd__decap_3 PHY_962 ();
 sky130_fd_sc_hd__decap_3 PHY_963 ();
 sky130_fd_sc_hd__decap_3 PHY_964 ();
 sky130_fd_sc_hd__decap_3 PHY_965 ();
 sky130_fd_sc_hd__decap_3 PHY_966 ();
 sky130_fd_sc_hd__decap_3 PHY_967 ();
 sky130_fd_sc_hd__decap_3 PHY_968 ();
 sky130_fd_sc_hd__decap_3 PHY_969 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_970 ();
 sky130_fd_sc_hd__decap_3 PHY_971 ();
 sky130_fd_sc_hd__decap_3 PHY_972 ();
 sky130_fd_sc_hd__decap_3 PHY_973 ();
 sky130_fd_sc_hd__decap_3 PHY_974 ();
 sky130_fd_sc_hd__decap_3 PHY_975 ();
 sky130_fd_sc_hd__decap_3 PHY_976 ();
 sky130_fd_sc_hd__decap_3 PHY_977 ();
 sky130_fd_sc_hd__decap_3 PHY_978 ();
 sky130_fd_sc_hd__decap_3 PHY_979 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_980 ();
 sky130_fd_sc_hd__decap_3 PHY_981 ();
 sky130_fd_sc_hd__decap_3 PHY_982 ();
 sky130_fd_sc_hd__decap_3 PHY_983 ();
 sky130_fd_sc_hd__decap_3 PHY_984 ();
 sky130_fd_sc_hd__decap_3 PHY_985 ();
 sky130_fd_sc_hd__decap_3 PHY_986 ();
 sky130_fd_sc_hd__decap_3 PHY_987 ();
 sky130_fd_sc_hd__decap_3 PHY_988 ();
 sky130_fd_sc_hd__decap_3 PHY_989 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_990 ();
 sky130_fd_sc_hd__decap_3 PHY_991 ();
 sky130_fd_sc_hd__decap_3 PHY_992 ();
 sky130_fd_sc_hd__decap_3 PHY_993 ();
 sky130_fd_sc_hd__decap_3 PHY_994 ();
 sky130_fd_sc_hd__decap_3 PHY_995 ();
 sky130_fd_sc_hd__decap_3 PHY_996 ();
 sky130_fd_sc_hd__decap_3 PHY_997 ();
 sky130_fd_sc_hd__decap_3 PHY_998 ();
 sky130_fd_sc_hd__decap_3 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__inv_2 _4098_ (.A(net144),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_2 _4099_ (.A(net16),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_2 _4100_ (.A(net15),
    .Y(_0561_));
 sky130_fd_sc_hd__inv_2 _4101_ (.A(net18),
    .Y(_0562_));
 sky130_fd_sc_hd__inv_2 _4102_ (.A(net17),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_2 _4103_ (.A(net31),
    .Y(_0564_));
 sky130_fd_sc_hd__inv_2 _4104_ (.A(net25),
    .Y(_0565_));
 sky130_fd_sc_hd__inv_2 _4105_ (.A(net67),
    .Y(_0566_));
 sky130_fd_sc_hd__inv_2 _4106_ (.A(net784),
    .Y(_0567_));
 sky130_fd_sc_hd__inv_2 _4107_ (.A(net631),
    .Y(_0568_));
 sky130_fd_sc_hd__clkinv_4 _4108_ (.A(\ann.temp[29] ),
    .Y(_0569_));
 sky130_fd_sc_hd__inv_2 _4109_ (.A(\ann.ReLU_out[9][28] ),
    .Y(_0570_));
 sky130_fd_sc_hd__clkinv_4 _4110_ (.A(\ann.temp[28] ),
    .Y(_0571_));
 sky130_fd_sc_hd__clkinv_4 _4111_ (.A(\ann.temp[27] ),
    .Y(_0572_));
 sky130_fd_sc_hd__inv_2 _4112_ (.A(net182),
    .Y(_0573_));
 sky130_fd_sc_hd__inv_2 _4113_ (.A(\ann.temp[25] ),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_2 _4114_ (.A(\ann.ReLU_out[9][24] ),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_2 _4115_ (.A(\ann.ReLU_out[9][23] ),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_2 _4116_ (.A(\ann.ReLU_out[9][22] ),
    .Y(_0577_));
 sky130_fd_sc_hd__inv_2 _4117_ (.A(\ann.temp[22] ),
    .Y(_0578_));
 sky130_fd_sc_hd__inv_4 _4118_ (.A(\ann.temp[21] ),
    .Y(_0579_));
 sky130_fd_sc_hd__inv_4 _4119_ (.A(\ann.temp[20] ),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_2 _4120_ (.A(\ann.ReLU_out[8][29] ),
    .Y(_0581_));
 sky130_fd_sc_hd__inv_2 _4121_ (.A(\ann.ReLU_out[8][26] ),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_2 _4122_ (.A(\ann.ReLU_out[8][25] ),
    .Y(_0583_));
 sky130_fd_sc_hd__inv_2 _4123_ (.A(\ann.ReLU_out[8][24] ),
    .Y(_0584_));
 sky130_fd_sc_hd__inv_2 _4124_ (.A(\ann.ReLU_out[8][23] ),
    .Y(_0585_));
 sky130_fd_sc_hd__inv_2 _4125_ (.A(\ann.ReLU_out[8][22] ),
    .Y(_0586_));
 sky130_fd_sc_hd__inv_2 _4126_ (.A(\ann.ReLU_out[8][21] ),
    .Y(_0587_));
 sky130_fd_sc_hd__inv_2 _4127_ (.A(\ann.ReLU_out[8][20] ),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_2 _4128_ (.A(\ann.ReLU_out[7][29] ),
    .Y(_0589_));
 sky130_fd_sc_hd__inv_2 _4129_ (.A(\ann.ReLU_out[7][26] ),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_2 _4130_ (.A(\ann.ReLU_out[7][25] ),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_2 _4131_ (.A(\ann.ReLU_out[7][24] ),
    .Y(_0592_));
 sky130_fd_sc_hd__inv_2 _4132_ (.A(\ann.ReLU_out[7][23] ),
    .Y(_0593_));
 sky130_fd_sc_hd__inv_2 _4133_ (.A(\ann.ReLU_out[7][22] ),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_2 _4134_ (.A(\ann.ReLU_out[7][21] ),
    .Y(_0595_));
 sky130_fd_sc_hd__inv_2 _4135_ (.A(\ann.ReLU_out[7][20] ),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _4136_ (.A(net321),
    .Y(_0597_));
 sky130_fd_sc_hd__inv_2 _4137_ (.A(\ann.ReLU_out[6][27] ),
    .Y(_0598_));
 sky130_fd_sc_hd__inv_2 _4138_ (.A(\ann.ReLU_out[6][26] ),
    .Y(_0599_));
 sky130_fd_sc_hd__inv_2 _4139_ (.A(\ann.ReLU_out[6][25] ),
    .Y(_0600_));
 sky130_fd_sc_hd__inv_2 _4140_ (.A(\ann.ReLU_out[6][24] ),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_2 _4141_ (.A(\ann.ReLU_out[6][23] ),
    .Y(_0602_));
 sky130_fd_sc_hd__inv_2 _4142_ (.A(\ann.ReLU_out[6][20] ),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _4143_ (.A(\ann.ReLU_out[5][29] ),
    .Y(_0604_));
 sky130_fd_sc_hd__inv_2 _4144_ (.A(\ann.ReLU_out[5][28] ),
    .Y(_0605_));
 sky130_fd_sc_hd__inv_2 _4145_ (.A(\ann.ReLU_out[5][27] ),
    .Y(_0606_));
 sky130_fd_sc_hd__inv_2 _4146_ (.A(\ann.ReLU_out[5][26] ),
    .Y(_0607_));
 sky130_fd_sc_hd__inv_2 _4147_ (.A(\ann.ReLU_out[5][25] ),
    .Y(_0608_));
 sky130_fd_sc_hd__inv_2 _4148_ (.A(\ann.ReLU_out[5][24] ),
    .Y(_0609_));
 sky130_fd_sc_hd__inv_2 _4149_ (.A(\ann.ReLU_out[5][23] ),
    .Y(_0610_));
 sky130_fd_sc_hd__inv_2 _4150_ (.A(\ann.ReLU_out[5][22] ),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _4151_ (.A(\ann.ReLU_out[4][29] ),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_2 _4152_ (.A(net674),
    .Y(_0613_));
 sky130_fd_sc_hd__inv_2 _4153_ (.A(\ann.ReLU_out[4][27] ),
    .Y(_0614_));
 sky130_fd_sc_hd__inv_2 _4154_ (.A(\ann.ReLU_out[4][26] ),
    .Y(_0615_));
 sky130_fd_sc_hd__inv_2 _4155_ (.A(\ann.ReLU_out[4][25] ),
    .Y(_0616_));
 sky130_fd_sc_hd__inv_2 _4156_ (.A(\ann.ReLU_out[4][24] ),
    .Y(_0617_));
 sky130_fd_sc_hd__inv_2 _4157_ (.A(\ann.ReLU_out[4][23] ),
    .Y(_0618_));
 sky130_fd_sc_hd__inv_2 _4158_ (.A(\ann.ReLU_out[4][22] ),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_2 _4159_ (.A(\ann.ReLU_out[3][25] ),
    .Y(_0620_));
 sky130_fd_sc_hd__inv_2 _4160_ (.A(\ann.ReLU_out[3][24] ),
    .Y(_0621_));
 sky130_fd_sc_hd__inv_2 _4161_ (.A(\ann.ReLU_out[3][23] ),
    .Y(_0622_));
 sky130_fd_sc_hd__inv_2 _4162_ (.A(\ann.ReLU_out[3][22] ),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _4163_ (.A(\ann.ReLU_out[2][29] ),
    .Y(_0624_));
 sky130_fd_sc_hd__inv_2 _4164_ (.A(net618),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_2 _4165_ (.A(\ann.ReLU_out[2][27] ),
    .Y(_0626_));
 sky130_fd_sc_hd__inv_2 _4166_ (.A(\ann.ReLU_out[2][26] ),
    .Y(_0627_));
 sky130_fd_sc_hd__inv_2 _4167_ (.A(\ann.ReLU_out[2][25] ),
    .Y(_0628_));
 sky130_fd_sc_hd__inv_2 _4168_ (.A(net437),
    .Y(_0629_));
 sky130_fd_sc_hd__inv_2 _4169_ (.A(\ann.ReLU_out[2][23] ),
    .Y(_0630_));
 sky130_fd_sc_hd__inv_2 _4170_ (.A(\ann.ReLU_out[2][22] ),
    .Y(_0631_));
 sky130_fd_sc_hd__inv_2 _4171_ (.A(\ann.ReLU_out[1][30] ),
    .Y(_0632_));
 sky130_fd_sc_hd__inv_2 _4172_ (.A(\ann.ReLU_out[1][27] ),
    .Y(_0633_));
 sky130_fd_sc_hd__inv_2 _4173_ (.A(\ann.ReLU_out[1][26] ),
    .Y(_0634_));
 sky130_fd_sc_hd__inv_2 _4174_ (.A(\ann.ReLU_out[1][25] ),
    .Y(_0635_));
 sky130_fd_sc_hd__inv_2 _4175_ (.A(net436),
    .Y(_0636_));
 sky130_fd_sc_hd__inv_2 _4176_ (.A(net432),
    .Y(_0637_));
 sky130_fd_sc_hd__inv_2 _4177_ (.A(\ann.ReLU_out[1][22] ),
    .Y(_0638_));
 sky130_fd_sc_hd__inv_2 _4178_ (.A(\ann.temp[19] ),
    .Y(_0639_));
 sky130_fd_sc_hd__inv_2 _4179_ (.A(net187),
    .Y(_0640_));
 sky130_fd_sc_hd__inv_2 _4180_ (.A(net456),
    .Y(_0641_));
 sky130_fd_sc_hd__inv_2 _4181_ (.A(net188),
    .Y(_0642_));
 sky130_fd_sc_hd__inv_2 _4182_ (.A(\ann.temp[16] ),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_2 _4183_ (.A(net410),
    .Y(_0644_));
 sky130_fd_sc_hd__inv_2 _4184_ (.A(\ann.ReLU_out[1][15] ),
    .Y(_0645_));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(\ann.temp[15] ),
    .Y(_0646_));
 sky130_fd_sc_hd__inv_2 _4186_ (.A(\ann.temp[14] ),
    .Y(_0647_));
 sky130_fd_sc_hd__inv_2 _4187_ (.A(\ann.temp[13] ),
    .Y(_0648_));
 sky130_fd_sc_hd__inv_2 _4188_ (.A(\ann.temp[12] ),
    .Y(_0649_));
 sky130_fd_sc_hd__inv_2 _4189_ (.A(\ann.temp[11] ),
    .Y(_0650_));
 sky130_fd_sc_hd__inv_2 _4190_ (.A(\ann.temp[10] ),
    .Y(_0651_));
 sky130_fd_sc_hd__inv_2 _4191_ (.A(\ann.temp[9] ),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _4192_ (.A(\ann.ReLU_out[1][8] ),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_2 _4193_ (.A(net333),
    .Y(_0654_));
 sky130_fd_sc_hd__inv_2 _4194_ (.A(net379),
    .Y(_0655_));
 sky130_fd_sc_hd__inv_2 _4195_ (.A(net329),
    .Y(_0656_));
 sky130_fd_sc_hd__inv_2 _4196_ (.A(\ann.temp[4] ),
    .Y(_0657_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(\ann.temp[3] ),
    .Y(_0658_));
 sky130_fd_sc_hd__inv_2 _4198_ (.A(\ann.temp[2] ),
    .Y(_0659_));
 sky130_fd_sc_hd__inv_2 _4199_ (.A(\ann.temp[1] ),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _4200_ (.A(\ann.temp[0] ),
    .Y(_0661_));
 sky130_fd_sc_hd__inv_2 _4201_ (.A(\ann.ReLU_out[2][18] ),
    .Y(_0662_));
 sky130_fd_sc_hd__inv_2 _4202_ (.A(\ann.ReLU_out[2][17] ),
    .Y(_0663_));
 sky130_fd_sc_hd__inv_2 _4203_ (.A(\ann.ReLU_out[2][15] ),
    .Y(_0664_));
 sky130_fd_sc_hd__inv_2 _4204_ (.A(\ann.ReLU_out[2][8] ),
    .Y(_0665_));
 sky130_fd_sc_hd__inv_2 _4205_ (.A(\ann.ReLU_out[3][18] ),
    .Y(_0666_));
 sky130_fd_sc_hd__inv_2 _4206_ (.A(\ann.ReLU_out[3][15] ),
    .Y(_0667_));
 sky130_fd_sc_hd__inv_2 _4207_ (.A(\ann.ReLU_out[3][8] ),
    .Y(_0668_));
 sky130_fd_sc_hd__inv_2 _4208_ (.A(net603),
    .Y(_0669_));
 sky130_fd_sc_hd__inv_2 _4209_ (.A(\ann.ReLU_out[4][17] ),
    .Y(_0670_));
 sky130_fd_sc_hd__inv_2 _4210_ (.A(\ann.ReLU_out[4][15] ),
    .Y(_0671_));
 sky130_fd_sc_hd__inv_2 _4211_ (.A(\ann.ReLU_out[4][8] ),
    .Y(_0672_));
 sky130_fd_sc_hd__inv_2 _4212_ (.A(\ann.ReLU_out[5][18] ),
    .Y(_0673_));
 sky130_fd_sc_hd__inv_2 _4213_ (.A(\ann.ReLU_out[5][17] ),
    .Y(_0674_));
 sky130_fd_sc_hd__inv_2 _4214_ (.A(\ann.ReLU_out[5][15] ),
    .Y(_0675_));
 sky130_fd_sc_hd__inv_2 _4215_ (.A(\ann.ReLU_out[5][8] ),
    .Y(_0676_));
 sky130_fd_sc_hd__inv_2 _4216_ (.A(\ann.ReLU_out[6][19] ),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_2 _4217_ (.A(\ann.ReLU_out[6][18] ),
    .Y(_0678_));
 sky130_fd_sc_hd__inv_2 _4218_ (.A(net335),
    .Y(_0679_));
 sky130_fd_sc_hd__inv_2 _4219_ (.A(net369),
    .Y(_0680_));
 sky130_fd_sc_hd__inv_2 _4220_ (.A(\ann.ReLU_out[6][15] ),
    .Y(_0681_));
 sky130_fd_sc_hd__inv_2 _4221_ (.A(\ann.ReLU_out[6][11] ),
    .Y(_0682_));
 sky130_fd_sc_hd__inv_2 _4222_ (.A(\ann.ReLU_out[6][10] ),
    .Y(_0683_));
 sky130_fd_sc_hd__inv_2 _4223_ (.A(\ann.ReLU_out[6][9] ),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _4224_ (.A(net337),
    .Y(_0685_));
 sky130_fd_sc_hd__inv_2 _4225_ (.A(\ann.ReLU_out[7][18] ),
    .Y(_0686_));
 sky130_fd_sc_hd__inv_2 _4226_ (.A(\ann.ReLU_out[7][17] ),
    .Y(_0687_));
 sky130_fd_sc_hd__inv_2 _4227_ (.A(\ann.ReLU_out[7][15] ),
    .Y(_0688_));
 sky130_fd_sc_hd__inv_2 _4228_ (.A(\ann.ReLU_out[7][11] ),
    .Y(_0689_));
 sky130_fd_sc_hd__inv_2 _4229_ (.A(\ann.ReLU_out[7][10] ),
    .Y(_0690_));
 sky130_fd_sc_hd__inv_2 _4230_ (.A(\ann.ReLU_out[7][9] ),
    .Y(_0691_));
 sky130_fd_sc_hd__inv_2 _4231_ (.A(\ann.ReLU_out[7][8] ),
    .Y(_0692_));
 sky130_fd_sc_hd__inv_2 _4232_ (.A(\ann.ReLU_out[8][18] ),
    .Y(_0693_));
 sky130_fd_sc_hd__inv_2 _4233_ (.A(\ann.ReLU_out[8][17] ),
    .Y(_0694_));
 sky130_fd_sc_hd__inv_2 _4234_ (.A(\ann.ReLU_out[8][15] ),
    .Y(_0695_));
 sky130_fd_sc_hd__inv_2 _4235_ (.A(\ann.ReLU_out[8][11] ),
    .Y(_0696_));
 sky130_fd_sc_hd__inv_2 _4236_ (.A(\ann.ReLU_out[8][10] ),
    .Y(_0697_));
 sky130_fd_sc_hd__inv_2 _4237_ (.A(\ann.ReLU_out[8][9] ),
    .Y(_0698_));
 sky130_fd_sc_hd__inv_2 _4238_ (.A(\ann.ReLU_out[8][8] ),
    .Y(_0699_));
 sky130_fd_sc_hd__inv_2 _4239_ (.A(\ann.ReLU_out[9][18] ),
    .Y(_0700_));
 sky130_fd_sc_hd__inv_2 _4240_ (.A(\ann.ReLU_out[9][17] ),
    .Y(_0701_));
 sky130_fd_sc_hd__inv_2 _4241_ (.A(\ann.ReLU_out[9][16] ),
    .Y(_0702_));
 sky130_fd_sc_hd__inv_2 _4242_ (.A(\ann.ReLU_out[9][15] ),
    .Y(_0703_));
 sky130_fd_sc_hd__inv_2 _4243_ (.A(\ann.ReLU_out[9][11] ),
    .Y(_0704_));
 sky130_fd_sc_hd__inv_2 _4244_ (.A(\ann.ReLU_out[9][10] ),
    .Y(_0705_));
 sky130_fd_sc_hd__inv_2 _4245_ (.A(\ann.ReLU_out[9][9] ),
    .Y(_0706_));
 sky130_fd_sc_hd__inv_2 _4246_ (.A(\ann.ReLU_out[9][8] ),
    .Y(_0707_));
 sky130_fd_sc_hd__and2b_1 _4247_ (.A_N(net731),
    .B(net402),
    .X(_0557_));
 sky130_fd_sc_hd__and2b_1 _4248_ (.A_N(net402),
    .B(net731),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_1 _4249_ (.A(net31),
    .B(net28),
    .Y(_0708_));
 sky130_fd_sc_hd__or2_2 _4250_ (.A(net31),
    .B(net28),
    .X(_0709_));
 sky130_fd_sc_hd__and3_1 _4251_ (.A(net145),
    .B(net180),
    .C(net207),
    .X(_0000_));
 sky130_fd_sc_hd__a22o_1 _4252_ (.A1(net143),
    .A2(net180),
    .B1(net178),
    .B2(net145),
    .X(_0710_));
 sky130_fd_sc_hd__and4_1 _4253_ (.A(net143),
    .B(net145),
    .C(net180),
    .D(net178),
    .X(_0711_));
 sky130_fd_sc_hd__and3b_1 _4254_ (.A_N(_0711_),
    .B(net207),
    .C(_0710_),
    .X(_0011_));
 sky130_fd_sc_hd__and4_1 _4255_ (.A(net140),
    .B(net143),
    .C(net180),
    .D(net178),
    .X(_0712_));
 sky130_fd_sc_hd__a22oi_1 _4256_ (.A1(net140),
    .A2(net180),
    .B1(net178),
    .B2(net143),
    .Y(_0713_));
 sky130_fd_sc_hd__nor2_1 _4257_ (.A(_0712_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__and3_1 _4258_ (.A(net145),
    .B(net177),
    .C(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__a21oi_1 _4259_ (.A1(net145),
    .A2(net177),
    .B1(_0714_),
    .Y(_0716_));
 sky130_fd_sc_hd__nor2_1 _4260_ (.A(_0715_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__and2_1 _4261_ (.A(_0711_),
    .B(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__o21ai_1 _4262_ (.A1(_0711_),
    .A2(_0717_),
    .B1(net207),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_1 _4263_ (.A(_0718_),
    .B(_0719_),
    .Y(_0022_));
 sky130_fd_sc_hd__nand2_1 _4264_ (.A(net145),
    .B(net175),
    .Y(_0720_));
 sky130_fd_sc_hd__nand2_1 _4265_ (.A(net143),
    .B(net177),
    .Y(_0721_));
 sky130_fd_sc_hd__and4_1 _4266_ (.A(net137),
    .B(net140),
    .C(net180),
    .D(net178),
    .X(_0722_));
 sky130_fd_sc_hd__a22o_1 _4267_ (.A1(net137),
    .A2(net180),
    .B1(net178),
    .B2(net140),
    .X(_0723_));
 sky130_fd_sc_hd__and2b_1 _4268_ (.A_N(_0722_),
    .B(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__xnor2_1 _4269_ (.A(_0721_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__o21ai_1 _4270_ (.A1(_0712_),
    .A2(_0715_),
    .B1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__or3_1 _4271_ (.A(_0712_),
    .B(_0715_),
    .C(_0725_),
    .X(_0727_));
 sky130_fd_sc_hd__and2_1 _4272_ (.A(_0726_),
    .B(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__nand2b_1 _4273_ (.A_N(_0720_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__xnor2_1 _4274_ (.A(_0720_),
    .B(_0728_),
    .Y(_0730_));
 sky130_fd_sc_hd__and2_1 _4275_ (.A(_0718_),
    .B(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__o21ai_1 _4276_ (.A1(_0718_),
    .A2(_0730_),
    .B1(net207),
    .Y(_0732_));
 sky130_fd_sc_hd__nor2_1 _4277_ (.A(_0731_),
    .B(_0732_),
    .Y(_0025_));
 sky130_fd_sc_hd__a22oi_1 _4278_ (.A1(net143),
    .A2(net175),
    .B1(net174),
    .B2(net145),
    .Y(_0733_));
 sky130_fd_sc_hd__and4_2 _4279_ (.A(net143),
    .B(net145),
    .C(net175),
    .D(net174),
    .X(_0734_));
 sky130_fd_sc_hd__nor2_1 _4280_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__a31o_1 _4281_ (.A1(net143),
    .A2(net177),
    .A3(_0723_),
    .B1(_0722_),
    .X(_0736_));
 sky130_fd_sc_hd__and2_1 _4282_ (.A(net140),
    .B(net177),
    .X(_0737_));
 sky130_fd_sc_hd__nand4_2 _4283_ (.A(net134),
    .B(net137),
    .C(net180),
    .D(net178),
    .Y(_0738_));
 sky130_fd_sc_hd__a22o_1 _4284_ (.A1(net134),
    .A2(net180),
    .B1(net178),
    .B2(net137),
    .X(_0739_));
 sky130_fd_sc_hd__nand3_1 _4285_ (.A(_0737_),
    .B(_0738_),
    .C(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__a21o_1 _4286_ (.A1(_0738_),
    .A2(_0739_),
    .B1(_0737_),
    .X(_0741_));
 sky130_fd_sc_hd__and3_1 _4287_ (.A(_0736_),
    .B(_0740_),
    .C(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__a21o_1 _4288_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0736_),
    .X(_0743_));
 sky130_fd_sc_hd__and2b_1 _4289_ (.A_N(_0742_),
    .B(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__xnor2_1 _4290_ (.A(_0735_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__a21o_2 _4291_ (.A1(_0726_),
    .A2(_0729_),
    .B1(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__nand3_1 _4292_ (.A(_0726_),
    .B(_0729_),
    .C(_0745_),
    .Y(_0747_));
 sky130_fd_sc_hd__a21o_1 _4293_ (.A1(_0746_),
    .A2(_0747_),
    .B1(_0731_),
    .X(_0748_));
 sky130_fd_sc_hd__nand3_2 _4294_ (.A(_0731_),
    .B(_0746_),
    .C(_0747_),
    .Y(_0749_));
 sky130_fd_sc_hd__and3_1 _4295_ (.A(net205),
    .B(_0748_),
    .C(_0749_),
    .X(_0026_));
 sky130_fd_sc_hd__a21o_1 _4296_ (.A1(_0735_),
    .A2(_0743_),
    .B1(_0742_),
    .X(_0750_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(net145),
    .B(net171),
    .Y(_0751_));
 sky130_fd_sc_hd__a22oi_1 _4298_ (.A1(net140),
    .A2(net175),
    .B1(net174),
    .B2(net143),
    .Y(_0752_));
 sky130_fd_sc_hd__and4_1 _4299_ (.A(net140),
    .B(net143),
    .C(net175),
    .D(net174),
    .X(_0753_));
 sky130_fd_sc_hd__nor2_1 _4300_ (.A(_0752_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__and3_1 _4301_ (.A(net145),
    .B(net171),
    .C(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__xnor2_1 _4302_ (.A(_0751_),
    .B(_0754_),
    .Y(_0756_));
 sky130_fd_sc_hd__a21bo_1 _4303_ (.A1(_0737_),
    .A2(_0739_),
    .B1_N(_0738_),
    .X(_0757_));
 sky130_fd_sc_hd__and2_1 _4304_ (.A(net137),
    .B(net177),
    .X(_0758_));
 sky130_fd_sc_hd__nand4_2 _4305_ (.A(net131),
    .B(net134),
    .C(net180),
    .D(net178),
    .Y(_0759_));
 sky130_fd_sc_hd__a22o_1 _4306_ (.A1(net131),
    .A2(net180),
    .B1(net178),
    .B2(net134),
    .X(_0760_));
 sky130_fd_sc_hd__nand3_1 _4307_ (.A(_0758_),
    .B(_0759_),
    .C(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__a21o_1 _4308_ (.A1(_0759_),
    .A2(_0760_),
    .B1(_0758_),
    .X(_0762_));
 sky130_fd_sc_hd__nand3_1 _4309_ (.A(_0757_),
    .B(_0761_),
    .C(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__a21o_1 _4310_ (.A1(_0761_),
    .A2(_0762_),
    .B1(_0757_),
    .X(_0764_));
 sky130_fd_sc_hd__nand3_1 _4311_ (.A(_0756_),
    .B(_0763_),
    .C(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__a21o_1 _4312_ (.A1(_0763_),
    .A2(_0764_),
    .B1(_0756_),
    .X(_0766_));
 sky130_fd_sc_hd__and3_1 _4313_ (.A(_0750_),
    .B(_0765_),
    .C(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__a21o_1 _4314_ (.A1(_0765_),
    .A2(_0766_),
    .B1(_0750_),
    .X(_0768_));
 sky130_fd_sc_hd__and2b_1 _4315_ (.A_N(_0767_),
    .B(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__xnor2_4 _4316_ (.A(_0734_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__xnor2_1 _4317_ (.A(_0746_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(_0749_),
    .B(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__o211a_1 _4319_ (.A1(_0749_),
    .A2(_0770_),
    .B1(_0772_),
    .C1(net208),
    .X(_0027_));
 sky130_fd_sc_hd__a21oi_1 _4320_ (.A1(_0734_),
    .A2(_0768_),
    .B1(_0767_),
    .Y(_0773_));
 sky130_fd_sc_hd__o211a_1 _4321_ (.A1(_0753_),
    .A2(_0755_),
    .B1(net145),
    .C1(net170),
    .X(_0774_));
 sky130_fd_sc_hd__a211oi_1 _4322_ (.A1(net145),
    .A2(net170),
    .B1(_0753_),
    .C1(_0755_),
    .Y(_0775_));
 sky130_fd_sc_hd__or2_1 _4323_ (.A(_0774_),
    .B(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__a21bo_1 _4324_ (.A1(_0756_),
    .A2(_0764_),
    .B1_N(_0763_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(net141),
    .B(net171),
    .Y(_0778_));
 sky130_fd_sc_hd__a22o_1 _4326_ (.A1(net137),
    .A2(net175),
    .B1(net174),
    .B2(net140),
    .X(_0779_));
 sky130_fd_sc_hd__and3_1 _4327_ (.A(net137),
    .B(net140),
    .C(net174),
    .X(_0780_));
 sky130_fd_sc_hd__a21bo_1 _4328_ (.A1(net175),
    .A2(_0780_),
    .B1_N(_0779_),
    .X(_0781_));
 sky130_fd_sc_hd__xor2_1 _4329_ (.A(_0778_),
    .B(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__a21bo_1 _4330_ (.A1(_0758_),
    .A2(_0760_),
    .B1_N(_0759_),
    .X(_0783_));
 sky130_fd_sc_hd__and2_1 _4331_ (.A(net134),
    .B(net177),
    .X(_0784_));
 sky130_fd_sc_hd__nand4_2 _4332_ (.A(net128),
    .B(net131),
    .C(net180),
    .D(net178),
    .Y(_0785_));
 sky130_fd_sc_hd__a22o_1 _4333_ (.A1(net128),
    .A2(net180),
    .B1(net178),
    .B2(net131),
    .X(_0786_));
 sky130_fd_sc_hd__nand3_1 _4334_ (.A(_0784_),
    .B(_0785_),
    .C(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__a21o_1 _4335_ (.A1(_0785_),
    .A2(_0786_),
    .B1(_0784_),
    .X(_0788_));
 sky130_fd_sc_hd__nand3_1 _4336_ (.A(_0783_),
    .B(_0787_),
    .C(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__a21o_1 _4337_ (.A1(_0787_),
    .A2(_0788_),
    .B1(_0783_),
    .X(_0790_));
 sky130_fd_sc_hd__nand3_1 _4338_ (.A(_0782_),
    .B(_0789_),
    .C(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__a21o_1 _4339_ (.A1(_0789_),
    .A2(_0790_),
    .B1(_0782_),
    .X(_0792_));
 sky130_fd_sc_hd__and3_2 _4340_ (.A(_0777_),
    .B(_0791_),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__a21oi_1 _4341_ (.A1(_0791_),
    .A2(_0792_),
    .B1(_0777_),
    .Y(_0794_));
 sky130_fd_sc_hd__nor3_2 _4342_ (.A(_0776_),
    .B(_0793_),
    .C(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__o21a_1 _4343_ (.A1(_0793_),
    .A2(_0794_),
    .B1(_0776_),
    .X(_0796_));
 sky130_fd_sc_hd__nor3_2 _4344_ (.A(_0773_),
    .B(_0795_),
    .C(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__o21a_1 _4345_ (.A1(_0795_),
    .A2(_0796_),
    .B1(_0773_),
    .X(_0798_));
 sky130_fd_sc_hd__nor4_2 _4346_ (.A(_0746_),
    .B(_0770_),
    .C(_0797_),
    .D(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__o22a_1 _4347_ (.A1(_0746_),
    .A2(_0770_),
    .B1(_0797_),
    .B2(_0798_),
    .X(_0800_));
 sky130_fd_sc_hd__o22a_1 _4348_ (.A1(_0749_),
    .A2(_0770_),
    .B1(_0799_),
    .B2(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__or4_2 _4349_ (.A(_0749_),
    .B(_0770_),
    .C(_0799_),
    .D(_0800_),
    .X(_0802_));
 sky130_fd_sc_hd__and3b_1 _4350_ (.A_N(_0801_),
    .B(_0802_),
    .C(net208),
    .X(_0028_));
 sky130_fd_sc_hd__and4_1 _4351_ (.A(net141),
    .B(net144),
    .C(net170),
    .D(net167),
    .X(_0803_));
 sky130_fd_sc_hd__a22oi_1 _4352_ (.A1(net141),
    .A2(net170),
    .B1(net167),
    .B2(net144),
    .Y(_0804_));
 sky130_fd_sc_hd__nor2_1 _4353_ (.A(_0803_),
    .B(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__a32o_1 _4354_ (.A1(net141),
    .A2(net171),
    .A3(_0779_),
    .B1(_0780_),
    .B2(net175),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_1 _4355_ (.A(_0805_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__or2_1 _4356_ (.A(_0805_),
    .B(_0806_),
    .X(_0808_));
 sky130_fd_sc_hd__and2_1 _4357_ (.A(_0807_),
    .B(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__a21bo_1 _4358_ (.A1(_0782_),
    .A2(_0790_),
    .B1_N(_0789_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_1 _4359_ (.A(net139),
    .B(net172),
    .Y(_0811_));
 sky130_fd_sc_hd__a22oi_1 _4360_ (.A1(net133),
    .A2(\ann.weight[3] ),
    .B1(net173),
    .B2(net135),
    .Y(_0812_));
 sky130_fd_sc_hd__and4_1 _4361_ (.A(net133),
    .B(net135),
    .C(\ann.weight[3] ),
    .D(net173),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_1 _4362_ (.A(_0812_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__xnor2_1 _4363_ (.A(_0811_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__a21bo_1 _4364_ (.A1(_0784_),
    .A2(_0786_),
    .B1_N(_0785_),
    .X(_0816_));
 sky130_fd_sc_hd__and2_1 _4365_ (.A(net131),
    .B(net177),
    .X(_0817_));
 sky130_fd_sc_hd__a22o_1 _4366_ (.A1(net126),
    .A2(net180),
    .B1(net178),
    .B2(net128),
    .X(_0818_));
 sky130_fd_sc_hd__nand4_1 _4367_ (.A(net126),
    .B(net128),
    .C(net180),
    .D(net179),
    .Y(_0819_));
 sky130_fd_sc_hd__nand3_1 _4368_ (.A(_0817_),
    .B(_0818_),
    .C(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a21o_1 _4369_ (.A1(_0818_),
    .A2(_0819_),
    .B1(_0817_),
    .X(_0821_));
 sky130_fd_sc_hd__nand3_1 _4370_ (.A(_0816_),
    .B(_0820_),
    .C(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21o_1 _4371_ (.A1(_0820_),
    .A2(_0821_),
    .B1(_0816_),
    .X(_0823_));
 sky130_fd_sc_hd__nand3_1 _4372_ (.A(_0815_),
    .B(_0822_),
    .C(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__a21o_1 _4373_ (.A1(_0822_),
    .A2(_0823_),
    .B1(_0815_),
    .X(_0825_));
 sky130_fd_sc_hd__nand3_2 _4374_ (.A(_0810_),
    .B(_0824_),
    .C(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_2 _4375_ (.A(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__a21o_1 _4376_ (.A1(_0824_),
    .A2(_0825_),
    .B1(_0810_),
    .X(_0828_));
 sky130_fd_sc_hd__and3_1 _4377_ (.A(_0809_),
    .B(_0826_),
    .C(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__nand3_2 _4378_ (.A(_0809_),
    .B(_0826_),
    .C(_0828_),
    .Y(_0830_));
 sky130_fd_sc_hd__a21o_1 _4379_ (.A1(_0826_),
    .A2(_0828_),
    .B1(_0809_),
    .X(_0831_));
 sky130_fd_sc_hd__o211ai_4 _4380_ (.A1(_0793_),
    .A2(_0795_),
    .B1(_0830_),
    .C1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__a211o_1 _4381_ (.A1(_0830_),
    .A2(_0831_),
    .B1(_0793_),
    .C1(_0795_),
    .X(_0833_));
 sky130_fd_sc_hd__nand3_2 _4382_ (.A(_0774_),
    .B(_0832_),
    .C(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21o_1 _4383_ (.A1(_0832_),
    .A2(_0833_),
    .B1(_0774_),
    .X(_0835_));
 sky130_fd_sc_hd__and2_2 _4384_ (.A(_0834_),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__or2_1 _4385_ (.A(_0797_),
    .B(_0799_),
    .X(_0837_));
 sky130_fd_sc_hd__xnor2_1 _4386_ (.A(_0836_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_1 _4387_ (.A(_0802_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__or2_1 _4388_ (.A(net195),
    .B(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__a21oi_1 _4389_ (.A1(_0802_),
    .A2(_0838_),
    .B1(_0840_),
    .Y(_0029_));
 sky130_fd_sc_hd__a22o_1 _4390_ (.A1(net139),
    .A2(net169),
    .B1(net166),
    .B2(net141),
    .X(_0841_));
 sky130_fd_sc_hd__nand4_1 _4391_ (.A(net139),
    .B(net141),
    .C(net169),
    .D(net166),
    .Y(_0842_));
 sky130_fd_sc_hd__a22oi_1 _4392_ (.A1(net144),
    .A2(net164),
    .B1(_0841_),
    .B2(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__and4_1 _4393_ (.A(net144),
    .B(net165),
    .C(_0841_),
    .D(_0842_),
    .X(_0844_));
 sky130_fd_sc_hd__or2_1 _4394_ (.A(_0843_),
    .B(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__a31o_1 _4395_ (.A1(net138),
    .A2(net172),
    .A3(_0814_),
    .B1(_0813_),
    .X(_0846_));
 sky130_fd_sc_hd__and2b_1 _4396_ (.A_N(_0845_),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__xnor2_1 _4397_ (.A(_0845_),
    .B(_0846_),
    .Y(_0848_));
 sky130_fd_sc_hd__and2_1 _4398_ (.A(_0803_),
    .B(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__xnor2_1 _4399_ (.A(_0803_),
    .B(_0848_),
    .Y(_0850_));
 sky130_fd_sc_hd__a21bo_1 _4400_ (.A1(_0815_),
    .A2(_0823_),
    .B1_N(_0822_),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _4401_ (.A(net136),
    .B(net171),
    .Y(_0852_));
 sky130_fd_sc_hd__a22oi_1 _4402_ (.A1(net130),
    .A2(net176),
    .B1(net173),
    .B2(net133),
    .Y(_0853_));
 sky130_fd_sc_hd__and4_1 _4403_ (.A(net130),
    .B(net133),
    .C(net176),
    .D(net173),
    .X(_0854_));
 sky130_fd_sc_hd__nor2_1 _4404_ (.A(_0853_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__xnor2_1 _4405_ (.A(_0852_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21bo_1 _4406_ (.A1(_0817_),
    .A2(_0818_),
    .B1_N(_0819_),
    .X(_0857_));
 sky130_fd_sc_hd__and2_1 _4407_ (.A(net128),
    .B(\ann.weight[2] ),
    .X(_0858_));
 sky130_fd_sc_hd__nand4_2 _4408_ (.A(net123),
    .B(net126),
    .C(net181),
    .D(net179),
    .Y(_0859_));
 sky130_fd_sc_hd__a22o_1 _4409_ (.A1(net123),
    .A2(net181),
    .B1(net179),
    .B2(net126),
    .X(_0860_));
 sky130_fd_sc_hd__nand3_1 _4410_ (.A(_0858_),
    .B(_0859_),
    .C(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__a21o_1 _4411_ (.A1(_0859_),
    .A2(_0860_),
    .B1(_0858_),
    .X(_0862_));
 sky130_fd_sc_hd__nand3_1 _4412_ (.A(_0857_),
    .B(_0861_),
    .C(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21o_1 _4413_ (.A1(_0861_),
    .A2(_0862_),
    .B1(_0857_),
    .X(_0864_));
 sky130_fd_sc_hd__nand3_1 _4414_ (.A(_0856_),
    .B(_0863_),
    .C(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__a21o_1 _4415_ (.A1(_0863_),
    .A2(_0864_),
    .B1(_0856_),
    .X(_0866_));
 sky130_fd_sc_hd__and3_1 _4416_ (.A(_0851_),
    .B(_0865_),
    .C(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__nand3_1 _4417_ (.A(_0851_),
    .B(_0865_),
    .C(_0866_),
    .Y(_0868_));
 sky130_fd_sc_hd__a21oi_1 _4418_ (.A1(_0865_),
    .A2(_0866_),
    .B1(_0851_),
    .Y(_0869_));
 sky130_fd_sc_hd__or3_2 _4419_ (.A(_0850_),
    .B(_0867_),
    .C(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__o21ai_2 _4420_ (.A1(_0867_),
    .A2(_0869_),
    .B1(_0850_),
    .Y(_0871_));
 sky130_fd_sc_hd__o211a_2 _4421_ (.A1(_0827_),
    .A2(_0829_),
    .B1(_0870_),
    .C1(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__a211oi_2 _4422_ (.A1(_0870_),
    .A2(_0871_),
    .B1(_0827_),
    .C1(_0829_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor3_4 _4423_ (.A(_0807_),
    .B(_0872_),
    .C(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__o21a_1 _4424_ (.A1(_0872_),
    .A2(_0873_),
    .B1(_0807_),
    .X(_0875_));
 sky130_fd_sc_hd__a211oi_4 _4425_ (.A1(_0832_),
    .A2(_0834_),
    .B1(_0874_),
    .C1(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__o211a_1 _4426_ (.A1(_0874_),
    .A2(_0875_),
    .B1(_0832_),
    .C1(_0834_),
    .X(_0877_));
 sky130_fd_sc_hd__o211ai_1 _4427_ (.A1(_0874_),
    .A2(_0875_),
    .B1(_0832_),
    .C1(_0834_),
    .Y(_0878_));
 sky130_fd_sc_hd__or4bb_2 _4428_ (.A(_0876_),
    .B(_0877_),
    .C_N(_0797_),
    .D_N(_0836_),
    .X(_0879_));
 sky130_fd_sc_hd__a2bb2o_1 _4429_ (.A1_N(_0876_),
    .A2_N(_0877_),
    .B1(_0797_),
    .B2(_0836_),
    .X(_0880_));
 sky130_fd_sc_hd__nand4_2 _4430_ (.A(_0799_),
    .B(_0836_),
    .C(_0879_),
    .D(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__a22o_1 _4431_ (.A1(_0799_),
    .A2(_0836_),
    .B1(_0879_),
    .B2(_0880_),
    .X(_0882_));
 sky130_fd_sc_hd__a21o_1 _4432_ (.A1(_0881_),
    .A2(_0882_),
    .B1(_0839_),
    .X(_0883_));
 sky130_fd_sc_hd__nand3_1 _4433_ (.A(_0839_),
    .B(_0881_),
    .C(_0882_),
    .Y(_0884_));
 sky130_fd_sc_hd__and3_1 _4434_ (.A(net208),
    .B(_0883_),
    .C(_0884_),
    .X(_0030_));
 sky130_fd_sc_hd__o211a_1 _4435_ (.A1(_0847_),
    .A2(_0849_),
    .B1(net144),
    .C1(net163),
    .X(_0885_));
 sky130_fd_sc_hd__a211oi_1 _4436_ (.A1(net144),
    .A2(net163),
    .B1(_0847_),
    .C1(_0849_),
    .Y(_0886_));
 sky130_fd_sc_hd__or2_1 _4437_ (.A(_0885_),
    .B(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__a41o_1 _4438_ (.A1(net138),
    .A2(net141),
    .A3(net168),
    .A4(\ann.weight[7] ),
    .B1(_0844_),
    .X(_0888_));
 sky130_fd_sc_hd__nand2_1 _4439_ (.A(net141),
    .B(net165),
    .Y(_0889_));
 sky130_fd_sc_hd__and4_1 _4440_ (.A(net135),
    .B(net139),
    .C(net169),
    .D(\ann.weight[7] ),
    .X(_0890_));
 sky130_fd_sc_hd__a22o_1 _4441_ (.A1(net135),
    .A2(net169),
    .B1(net167),
    .B2(net139),
    .X(_0891_));
 sky130_fd_sc_hd__and2b_1 _4442_ (.A_N(_0890_),
    .B(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__xnor2_1 _4443_ (.A(_0889_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__o21ba_1 _4444_ (.A1(_0852_),
    .A2(_0853_),
    .B1_N(_0854_),
    .X(_0894_));
 sky130_fd_sc_hd__and2b_1 _4445_ (.A_N(_0894_),
    .B(_0893_),
    .X(_0895_));
 sky130_fd_sc_hd__xnor2_1 _4446_ (.A(_0893_),
    .B(_0894_),
    .Y(_0896_));
 sky130_fd_sc_hd__and2_1 _4447_ (.A(_0888_),
    .B(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__xor2_1 _4448_ (.A(_0888_),
    .B(_0896_),
    .X(_0898_));
 sky130_fd_sc_hd__a21bo_1 _4449_ (.A1(_0856_),
    .A2(_0864_),
    .B1_N(_0863_),
    .X(_0899_));
 sky130_fd_sc_hd__nand2_1 _4450_ (.A(net133),
    .B(net172),
    .Y(_0900_));
 sky130_fd_sc_hd__a22oi_2 _4451_ (.A1(net127),
    .A2(net176),
    .B1(net173),
    .B2(net129),
    .Y(_0901_));
 sky130_fd_sc_hd__and4_1 _4452_ (.A(net127),
    .B(net129),
    .C(net176),
    .D(net173),
    .X(_0902_));
 sky130_fd_sc_hd__nor2_1 _4453_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__xnor2_2 _4454_ (.A(_0900_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__a21bo_1 _4455_ (.A1(_0858_),
    .A2(_0860_),
    .B1_N(_0859_),
    .X(_0905_));
 sky130_fd_sc_hd__and2_1 _4456_ (.A(\ann.in_ff[2][7] ),
    .B(net177),
    .X(_0906_));
 sky130_fd_sc_hd__a22o_1 _4457_ (.A1(net120),
    .A2(net181),
    .B1(net179),
    .B2(\ann.in_ff[2][8] ),
    .X(_0907_));
 sky130_fd_sc_hd__nand4_2 _4458_ (.A(net120),
    .B(\ann.in_ff[2][8] ),
    .C(net181),
    .D(net179),
    .Y(_0908_));
 sky130_fd_sc_hd__nand3_1 _4459_ (.A(_0906_),
    .B(_0907_),
    .C(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21o_1 _4460_ (.A1(_0907_),
    .A2(_0908_),
    .B1(_0906_),
    .X(_0910_));
 sky130_fd_sc_hd__nand3_1 _4461_ (.A(_0905_),
    .B(_0909_),
    .C(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__a21o_1 _4462_ (.A1(_0909_),
    .A2(_0910_),
    .B1(_0905_),
    .X(_0912_));
 sky130_fd_sc_hd__nand3_1 _4463_ (.A(_0904_),
    .B(_0911_),
    .C(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__a21o_1 _4464_ (.A1(_0911_),
    .A2(_0912_),
    .B1(_0904_),
    .X(_0914_));
 sky130_fd_sc_hd__nand3_2 _4465_ (.A(_0899_),
    .B(_0913_),
    .C(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__a21o_1 _4466_ (.A1(_0913_),
    .A2(_0914_),
    .B1(_0899_),
    .X(_0916_));
 sky130_fd_sc_hd__and3_1 _4467_ (.A(_0898_),
    .B(_0915_),
    .C(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__nand3_1 _4468_ (.A(_0898_),
    .B(_0915_),
    .C(_0916_),
    .Y(_0918_));
 sky130_fd_sc_hd__a21oi_1 _4469_ (.A1(_0915_),
    .A2(_0916_),
    .B1(_0898_),
    .Y(_0919_));
 sky130_fd_sc_hd__a211oi_1 _4470_ (.A1(_0868_),
    .A2(_0870_),
    .B1(_0917_),
    .C1(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__a211o_1 _4471_ (.A1(_0868_),
    .A2(_0870_),
    .B1(_0917_),
    .C1(_0919_),
    .X(_0921_));
 sky130_fd_sc_hd__o211a_1 _4472_ (.A1(_0917_),
    .A2(_0919_),
    .B1(_0868_),
    .C1(_0870_),
    .X(_0922_));
 sky130_fd_sc_hd__or3_2 _4473_ (.A(_0887_),
    .B(_0920_),
    .C(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__o21ai_1 _4474_ (.A1(_0920_),
    .A2(_0922_),
    .B1(_0887_),
    .Y(_0924_));
 sky130_fd_sc_hd__o211a_1 _4475_ (.A1(_0872_),
    .A2(_0874_),
    .B1(_0923_),
    .C1(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__a211o_1 _4476_ (.A1(_0923_),
    .A2(_0924_),
    .B1(_0872_),
    .C1(_0874_),
    .X(_0926_));
 sky130_fd_sc_hd__and2b_1 _4477_ (.A_N(_0925_),
    .B(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__a31o_1 _4478_ (.A1(_0797_),
    .A2(_0836_),
    .A3(_0878_),
    .B1(_0876_),
    .X(_0928_));
 sky130_fd_sc_hd__xor2_1 _4479_ (.A(_0927_),
    .B(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__nand2b_1 _4480_ (.A_N(_0881_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2b_1 _4481_ (.A_N(_0929_),
    .B(_0881_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_0930_),
    .B(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__and2b_1 _4483_ (.A_N(_0884_),
    .B(_0929_),
    .X(_0933_));
 sky130_fd_sc_hd__a211oi_1 _4484_ (.A1(_0884_),
    .A2(_0932_),
    .B1(_0933_),
    .C1(net195),
    .Y(_0031_));
 sky130_fd_sc_hd__nand2b_1 _4485_ (.A_N(_0879_),
    .B(_0927_),
    .Y(_0934_));
 sky130_fd_sc_hd__a22oi_1 _4486_ (.A1(net141),
    .A2(net162),
    .B1(net158),
    .B2(net144),
    .Y(_0935_));
 sky130_fd_sc_hd__and4_1 _4487_ (.A(net141),
    .B(net144),
    .C(net161),
    .D(net158),
    .X(_0936_));
 sky130_fd_sc_hd__nor2_1 _4488_ (.A(_0935_),
    .B(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__o21ai_2 _4489_ (.A1(_0895_),
    .A2(_0897_),
    .B1(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__or3_1 _4490_ (.A(_0895_),
    .B(_0897_),
    .C(_0937_),
    .X(_0939_));
 sky130_fd_sc_hd__and2_1 _4491_ (.A(_0938_),
    .B(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__a31o_1 _4492_ (.A1(net142),
    .A2(net164),
    .A3(_0891_),
    .B1(_0890_),
    .X(_0941_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(net138),
    .B(net165),
    .Y(_0942_));
 sky130_fd_sc_hd__a22o_1 _4494_ (.A1(net132),
    .A2(net168),
    .B1(net167),
    .B2(net136),
    .X(_0943_));
 sky130_fd_sc_hd__and3_1 _4495_ (.A(net132),
    .B(net136),
    .C(net167),
    .X(_0944_));
 sky130_fd_sc_hd__a21bo_1 _4496_ (.A1(net168),
    .A2(_0944_),
    .B1_N(_0943_),
    .X(_0945_));
 sky130_fd_sc_hd__xor2_1 _4497_ (.A(_0942_),
    .B(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__o21ba_1 _4498_ (.A1(_0900_),
    .A2(_0901_),
    .B1_N(_0902_),
    .X(_0947_));
 sky130_fd_sc_hd__nand2b_1 _4499_ (.A_N(_0947_),
    .B(_0946_),
    .Y(_0948_));
 sky130_fd_sc_hd__xnor2_1 _4500_ (.A(_0946_),
    .B(_0947_),
    .Y(_0949_));
 sky130_fd_sc_hd__nand2_1 _4501_ (.A(_0941_),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__xor2_1 _4502_ (.A(_0941_),
    .B(_0949_),
    .X(_0951_));
 sky130_fd_sc_hd__a21bo_1 _4503_ (.A1(_0904_),
    .A2(_0912_),
    .B1_N(_0911_),
    .X(_0952_));
 sky130_fd_sc_hd__nand2_1 _4504_ (.A(net129),
    .B(net171),
    .Y(_0953_));
 sky130_fd_sc_hd__a22o_1 _4505_ (.A1(net125),
    .A2(net176),
    .B1(net173),
    .B2(net127),
    .X(_0954_));
 sky130_fd_sc_hd__and3_1 _4506_ (.A(net126),
    .B(net127),
    .C(net173),
    .X(_0955_));
 sky130_fd_sc_hd__a21bo_1 _4507_ (.A1(net176),
    .A2(_0955_),
    .B1_N(_0954_),
    .X(_0956_));
 sky130_fd_sc_hd__xor2_2 _4508_ (.A(_0953_),
    .B(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__a21bo_1 _4509_ (.A1(_0906_),
    .A2(_0907_),
    .B1_N(_0908_),
    .X(_0958_));
 sky130_fd_sc_hd__and2_1 _4510_ (.A(\ann.in_ff[2][8] ),
    .B(\ann.weight[2] ),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _4511_ (.A1(net118),
    .A2(\ann.weight[0] ),
    .B1(net179),
    .B2(net120),
    .X(_0960_));
 sky130_fd_sc_hd__nand4_1 _4512_ (.A(net118),
    .B(net120),
    .C(net181),
    .D(net179),
    .Y(_0961_));
 sky130_fd_sc_hd__nand3_1 _4513_ (.A(_0959_),
    .B(_0960_),
    .C(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__a21o_1 _4514_ (.A1(_0960_),
    .A2(_0961_),
    .B1(_0959_),
    .X(_0963_));
 sky130_fd_sc_hd__nand3_1 _4515_ (.A(_0958_),
    .B(_0962_),
    .C(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__a21o_1 _4516_ (.A1(_0962_),
    .A2(_0963_),
    .B1(_0958_),
    .X(_0965_));
 sky130_fd_sc_hd__nand3_2 _4517_ (.A(_0957_),
    .B(_0964_),
    .C(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__a21o_1 _4518_ (.A1(_0964_),
    .A2(_0965_),
    .B1(_0957_),
    .X(_0967_));
 sky130_fd_sc_hd__nand3_4 _4519_ (.A(_0952_),
    .B(_0966_),
    .C(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__a21o_1 _4520_ (.A1(_0966_),
    .A2(_0967_),
    .B1(_0952_),
    .X(_0969_));
 sky130_fd_sc_hd__and3_1 _4521_ (.A(_0951_),
    .B(_0968_),
    .C(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__nand3_2 _4522_ (.A(_0951_),
    .B(_0968_),
    .C(_0969_),
    .Y(_0971_));
 sky130_fd_sc_hd__a21oi_1 _4523_ (.A1(_0968_),
    .A2(_0969_),
    .B1(_0951_),
    .Y(_0972_));
 sky130_fd_sc_hd__a211o_2 _4524_ (.A1(_0915_),
    .A2(_0918_),
    .B1(_0970_),
    .C1(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__o211ai_2 _4525_ (.A1(_0970_),
    .A2(_0972_),
    .B1(_0915_),
    .C1(_0918_),
    .Y(_0974_));
 sky130_fd_sc_hd__and3_1 _4526_ (.A(_0940_),
    .B(_0973_),
    .C(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__nand3_1 _4527_ (.A(_0940_),
    .B(_0973_),
    .C(_0974_),
    .Y(_0976_));
 sky130_fd_sc_hd__a21oi_1 _4528_ (.A1(_0973_),
    .A2(_0974_),
    .B1(_0940_),
    .Y(_0977_));
 sky130_fd_sc_hd__a211o_2 _4529_ (.A1(_0921_),
    .A2(_0923_),
    .B1(_0975_),
    .C1(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__o211ai_2 _4530_ (.A1(_0975_),
    .A2(_0977_),
    .B1(_0921_),
    .C1(_0923_),
    .Y(_0979_));
 sky130_fd_sc_hd__and3_1 _4531_ (.A(_0885_),
    .B(_0978_),
    .C(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__nand3_1 _4532_ (.A(_0885_),
    .B(_0978_),
    .C(_0979_),
    .Y(_0981_));
 sky130_fd_sc_hd__a21oi_1 _4533_ (.A1(_0978_),
    .A2(_0979_),
    .B1(_0885_),
    .Y(_0982_));
 sky130_fd_sc_hd__nor2_1 _4534_ (.A(_0980_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__a21o_1 _4535_ (.A1(_0876_),
    .A2(_0926_),
    .B1(_0925_),
    .X(_0984_));
 sky130_fd_sc_hd__or3_1 _4536_ (.A(_0980_),
    .B(_0982_),
    .C(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__o21ai_1 _4537_ (.A1(_0980_),
    .A2(_0982_),
    .B1(_0984_),
    .Y(_0986_));
 sky130_fd_sc_hd__a21oi_2 _4538_ (.A1(_0985_),
    .A2(_0986_),
    .B1(_0934_),
    .Y(_0987_));
 sky130_fd_sc_hd__and3_1 _4539_ (.A(_0934_),
    .B(_0985_),
    .C(_0986_),
    .X(_0988_));
 sky130_fd_sc_hd__or3_1 _4540_ (.A(_0930_),
    .B(_0987_),
    .C(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__o21ai_2 _4541_ (.A1(_0987_),
    .A2(_0988_),
    .B1(_0930_),
    .Y(_0990_));
 sky130_fd_sc_hd__a21oi_1 _4542_ (.A1(_0989_),
    .A2(_0990_),
    .B1(_0933_),
    .Y(_0991_));
 sky130_fd_sc_hd__a31o_1 _4543_ (.A1(_0933_),
    .A2(_0989_),
    .A3(_0990_),
    .B1(net195),
    .X(_0992_));
 sky130_fd_sc_hd__nor2_1 _4544_ (.A(_0991_),
    .B(_0992_),
    .Y(_0001_));
 sky130_fd_sc_hd__a21bo_1 _4545_ (.A1(_0933_),
    .A2(_0990_),
    .B1_N(_0989_),
    .X(_0993_));
 sky130_fd_sc_hd__a22oi_1 _4546_ (.A1(net138),
    .A2(net161),
    .B1(net158),
    .B2(net141),
    .Y(_0994_));
 sky130_fd_sc_hd__and4_1 _4547_ (.A(net139),
    .B(net141),
    .C(net161),
    .D(net158),
    .X(_0995_));
 sky130_fd_sc_hd__and4bb_1 _4548_ (.A_N(_0994_),
    .B_N(_0995_),
    .C(net144),
    .D(net156),
    .X(_0996_));
 sky130_fd_sc_hd__o2bb2a_1 _4549_ (.A1_N(net144),
    .A2_N(net156),
    .B1(_0994_),
    .B2(_0995_),
    .X(_0997_));
 sky130_fd_sc_hd__nor2_1 _4550_ (.A(_0996_),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__and2_1 _4551_ (.A(_0936_),
    .B(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__xnor2_1 _4552_ (.A(_0936_),
    .B(_0998_),
    .Y(_1000_));
 sky130_fd_sc_hd__a21oi_1 _4553_ (.A1(_0948_),
    .A2(_0950_),
    .B1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__inv_2 _4554_ (.A(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__and3_1 _4555_ (.A(_0948_),
    .B(_0950_),
    .C(_1000_),
    .X(_1003_));
 sky130_fd_sc_hd__or2_1 _4556_ (.A(_1001_),
    .B(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__a32o_1 _4557_ (.A1(net139),
    .A2(net165),
    .A3(_0943_),
    .B1(_0944_),
    .B2(net168),
    .X(_1005_));
 sky130_fd_sc_hd__a22o_1 _4558_ (.A1(net129),
    .A2(net169),
    .B1(net166),
    .B2(net133),
    .X(_1006_));
 sky130_fd_sc_hd__and4_1 _4559_ (.A(net130),
    .B(net132),
    .C(net169),
    .D(net166),
    .X(_1007_));
 sky130_fd_sc_hd__nand4_1 _4560_ (.A(net130),
    .B(net133),
    .C(net168),
    .D(\ann.weight[7] ),
    .Y(_1008_));
 sky130_fd_sc_hd__and4_1 _4561_ (.A(net136),
    .B(net165),
    .C(_1006_),
    .D(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__a22o_1 _4562_ (.A1(net136),
    .A2(net164),
    .B1(_1006_),
    .B2(_1008_),
    .X(_1010_));
 sky130_fd_sc_hd__nand2b_1 _4563_ (.A_N(_1009_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__a32o_1 _4564_ (.A1(net130),
    .A2(net171),
    .A3(_0954_),
    .B1(_0955_),
    .B2(net176),
    .X(_1012_));
 sky130_fd_sc_hd__and2b_1 _4565_ (.A_N(_1011_),
    .B(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__xnor2_2 _4566_ (.A(_1011_),
    .B(_1012_),
    .Y(_1014_));
 sky130_fd_sc_hd__xor2_2 _4567_ (.A(_1005_),
    .B(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a21bo_1 _4568_ (.A1(_0957_),
    .A2(_0965_),
    .B1_N(_0964_),
    .X(_1016_));
 sky130_fd_sc_hd__nand2_1 _4569_ (.A(\ann.in_ff[2][6] ),
    .B(net171),
    .Y(_1017_));
 sky130_fd_sc_hd__a22oi_2 _4570_ (.A1(\ann.in_ff[2][8] ),
    .A2(\ann.weight[3] ),
    .B1(\ann.weight[4] ),
    .B2(\ann.in_ff[2][7] ),
    .Y(_1018_));
 sky130_fd_sc_hd__and4_1 _4571_ (.A(net123),
    .B(net125),
    .C(net176),
    .D(\ann.weight[4] ),
    .X(_1019_));
 sky130_fd_sc_hd__nor2_1 _4572_ (.A(_1018_),
    .B(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__xnor2_2 _4573_ (.A(_1017_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__a21bo_1 _4574_ (.A1(_0959_),
    .A2(_0960_),
    .B1_N(_0961_),
    .X(_1022_));
 sky130_fd_sc_hd__and2_1 _4575_ (.A(net120),
    .B(\ann.weight[2] ),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _4576_ (.A1(net114),
    .A2(\ann.weight[0] ),
    .B1(net179),
    .B2(net118),
    .X(_1024_));
 sky130_fd_sc_hd__nand4_1 _4577_ (.A(net114),
    .B(net117),
    .C(net181),
    .D(net179),
    .Y(_1025_));
 sky130_fd_sc_hd__nand3_1 _4578_ (.A(_1023_),
    .B(_1024_),
    .C(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__a21o_1 _4579_ (.A1(_1024_),
    .A2(_1025_),
    .B1(_1023_),
    .X(_1027_));
 sky130_fd_sc_hd__nand3_1 _4580_ (.A(_1022_),
    .B(_1026_),
    .C(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__a21o_1 _4581_ (.A1(_1026_),
    .A2(_1027_),
    .B1(_1022_),
    .X(_1029_));
 sky130_fd_sc_hd__nand3_2 _4582_ (.A(_1021_),
    .B(_1028_),
    .C(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__a21o_1 _4583_ (.A1(_1028_),
    .A2(_1029_),
    .B1(_1021_),
    .X(_1031_));
 sky130_fd_sc_hd__nand3_4 _4584_ (.A(_1016_),
    .B(_1030_),
    .C(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__a21o_1 _4585_ (.A1(_1030_),
    .A2(_1031_),
    .B1(_1016_),
    .X(_1033_));
 sky130_fd_sc_hd__and3_1 _4586_ (.A(_1015_),
    .B(_1032_),
    .C(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__nand3_2 _4587_ (.A(_1015_),
    .B(_1032_),
    .C(_1033_),
    .Y(_1035_));
 sky130_fd_sc_hd__a21oi_2 _4588_ (.A1(_1032_),
    .A2(_1033_),
    .B1(_1015_),
    .Y(_1036_));
 sky130_fd_sc_hd__a211oi_4 _4589_ (.A1(_0968_),
    .A2(_0971_),
    .B1(_1034_),
    .C1(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__o211a_1 _4590_ (.A1(_1034_),
    .A2(_1036_),
    .B1(_0968_),
    .C1(_0971_),
    .X(_1038_));
 sky130_fd_sc_hd__nor3_2 _4591_ (.A(_1004_),
    .B(_1037_),
    .C(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__o21a_1 _4592_ (.A1(_1037_),
    .A2(_1038_),
    .B1(_1004_),
    .X(_1040_));
 sky130_fd_sc_hd__a211oi_2 _4593_ (.A1(_0973_),
    .A2(_0976_),
    .B1(_1039_),
    .C1(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__o211a_1 _4594_ (.A1(_1039_),
    .A2(_1040_),
    .B1(_0973_),
    .C1(_0976_),
    .X(_1042_));
 sky130_fd_sc_hd__nor3_2 _4595_ (.A(_0938_),
    .B(_1041_),
    .C(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__o21a_1 _4596_ (.A1(_1041_),
    .A2(_1042_),
    .B1(_0938_),
    .X(_1044_));
 sky130_fd_sc_hd__a211oi_1 _4597_ (.A1(_0978_),
    .A2(_0981_),
    .B1(_1043_),
    .C1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a211o_1 _4598_ (.A1(_0978_),
    .A2(_0981_),
    .B1(_1043_),
    .C1(_1044_),
    .X(_1046_));
 sky130_fd_sc_hd__o211ai_2 _4599_ (.A1(_1043_),
    .A2(_1044_),
    .B1(_0978_),
    .C1(_0981_),
    .Y(_1047_));
 sky130_fd_sc_hd__nand4_2 _4600_ (.A(_0925_),
    .B(_0983_),
    .C(_1046_),
    .D(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__a22o_1 _4601_ (.A1(_0925_),
    .A2(_0983_),
    .B1(_1046_),
    .B2(_1047_),
    .X(_1049_));
 sky130_fd_sc_hd__nand3_1 _4602_ (.A(_0876_),
    .B(_0927_),
    .C(_0983_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand3b_2 _4603_ (.A_N(_1050_),
    .B(_1049_),
    .C(_1048_),
    .Y(_1051_));
 sky130_fd_sc_hd__a21bo_1 _4604_ (.A1(_1048_),
    .A2(_1049_),
    .B1_N(_1050_),
    .X(_1052_));
 sky130_fd_sc_hd__nand2_1 _4605_ (.A(_1051_),
    .B(_1052_),
    .Y(_1053_));
 sky130_fd_sc_hd__xor2_1 _4606_ (.A(_0993_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nand2_1 _4607_ (.A(_0987_),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__or2_1 _4608_ (.A(_0987_),
    .B(_1054_),
    .X(_1056_));
 sky130_fd_sc_hd__a21oi_1 _4609_ (.A1(_1055_),
    .A2(_1056_),
    .B1(net195),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(net145),
    .B(net154),
    .Y(_1057_));
 sky130_fd_sc_hd__or2_1 _4611_ (.A(_0995_),
    .B(_0996_),
    .X(_1058_));
 sky130_fd_sc_hd__a22oi_1 _4612_ (.A1(net136),
    .A2(net162),
    .B1(net159),
    .B2(net139),
    .Y(_1059_));
 sky130_fd_sc_hd__and4_1 _4613_ (.A(net136),
    .B(net139),
    .C(net162),
    .D(net159),
    .X(_1060_));
 sky130_fd_sc_hd__and4bb_1 _4614_ (.A_N(_1059_),
    .B_N(_1060_),
    .C(net141),
    .D(net156),
    .X(_1061_));
 sky130_fd_sc_hd__o2bb2a_1 _4615_ (.A1_N(net141),
    .A2_N(net156),
    .B1(_1059_),
    .B2(_1060_),
    .X(_1062_));
 sky130_fd_sc_hd__nor2_1 _4616_ (.A(_1061_),
    .B(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__nand2_1 _4617_ (.A(_1058_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__xor2_1 _4618_ (.A(_1058_),
    .B(_1063_),
    .X(_1065_));
 sky130_fd_sc_hd__nand2b_1 _4619_ (.A_N(_1057_),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__xnor2_1 _4620_ (.A(_1057_),
    .B(_1065_),
    .Y(_1067_));
 sky130_fd_sc_hd__a21oi_1 _4621_ (.A1(_1005_),
    .A2(_1014_),
    .B1(_1013_),
    .Y(_1068_));
 sky130_fd_sc_hd__and2b_1 _4622_ (.A_N(_1068_),
    .B(_1067_),
    .X(_1069_));
 sky130_fd_sc_hd__xnor2_1 _4623_ (.A(_1067_),
    .B(_1068_),
    .Y(_1070_));
 sky130_fd_sc_hd__xnor2_1 _4624_ (.A(_0999_),
    .B(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__nor2_1 _4625_ (.A(_1007_),
    .B(_1009_),
    .Y(_1072_));
 sky130_fd_sc_hd__a22oi_1 _4626_ (.A1(\ann.in_ff[2][6] ),
    .A2(net169),
    .B1(net166),
    .B2(net130),
    .Y(_1073_));
 sky130_fd_sc_hd__and4_1 _4627_ (.A(\ann.in_ff[2][6] ),
    .B(net130),
    .C(net169),
    .D(net166),
    .X(_1074_));
 sky130_fd_sc_hd__and4bb_1 _4628_ (.A_N(_1073_),
    .B_N(_1074_),
    .C(net133),
    .D(net164),
    .X(_1075_));
 sky130_fd_sc_hd__o2bb2a_1 _4629_ (.A1_N(net133),
    .A2_N(net164),
    .B1(_1073_),
    .B2(_1074_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_1 _4630_ (.A(_1075_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__o21ba_1 _4631_ (.A1(_1017_),
    .A2(_1018_),
    .B1_N(_1019_),
    .X(_1078_));
 sky130_fd_sc_hd__or3_1 _4632_ (.A(_1075_),
    .B(_1076_),
    .C(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__xnor2_1 _4633_ (.A(_1077_),
    .B(_1078_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2b_1 _4634_ (.A_N(_1072_),
    .B(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__xnor2_1 _4635_ (.A(_1072_),
    .B(_1080_),
    .Y(_1082_));
 sky130_fd_sc_hd__a21bo_1 _4636_ (.A1(_1021_),
    .A2(_1029_),
    .B1_N(_1028_),
    .X(_1083_));
 sky130_fd_sc_hd__nand2_1 _4637_ (.A(\ann.in_ff[2][7] ),
    .B(net172),
    .Y(_1084_));
 sky130_fd_sc_hd__a22oi_2 _4638_ (.A1(net121),
    .A2(net176),
    .B1(net173),
    .B2(net124),
    .Y(_1085_));
 sky130_fd_sc_hd__and4_1 _4639_ (.A(net121),
    .B(net124),
    .C(net176),
    .D(net173),
    .X(_1086_));
 sky130_fd_sc_hd__nor2_1 _4640_ (.A(_1085_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__xnor2_2 _4641_ (.A(_1084_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__a21bo_1 _4642_ (.A1(_1023_),
    .A2(_1024_),
    .B1_N(_1025_),
    .X(_1089_));
 sky130_fd_sc_hd__and2_1 _4643_ (.A(net117),
    .B(net177),
    .X(_1090_));
 sky130_fd_sc_hd__a22o_1 _4644_ (.A1(net111),
    .A2(\ann.weight[0] ),
    .B1(\ann.weight[1] ),
    .B2(net114),
    .X(_1091_));
 sky130_fd_sc_hd__nand4_1 _4645_ (.A(net111),
    .B(net114),
    .C(net181),
    .D(\ann.weight[1] ),
    .Y(_1092_));
 sky130_fd_sc_hd__nand3_1 _4646_ (.A(_1090_),
    .B(_1091_),
    .C(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__a21o_1 _4647_ (.A1(_1091_),
    .A2(_1092_),
    .B1(_1090_),
    .X(_1094_));
 sky130_fd_sc_hd__nand3_1 _4648_ (.A(_1089_),
    .B(_1093_),
    .C(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__a21o_1 _4649_ (.A1(_1093_),
    .A2(_1094_),
    .B1(_1089_),
    .X(_1096_));
 sky130_fd_sc_hd__nand3_2 _4650_ (.A(_1088_),
    .B(_1095_),
    .C(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__a21o_1 _4651_ (.A1(_1095_),
    .A2(_1096_),
    .B1(_1088_),
    .X(_1098_));
 sky130_fd_sc_hd__nand3_4 _4652_ (.A(_1083_),
    .B(_1097_),
    .C(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__a21o_1 _4653_ (.A1(_1097_),
    .A2(_1098_),
    .B1(_1083_),
    .X(_1100_));
 sky130_fd_sc_hd__and3_1 _4654_ (.A(_1082_),
    .B(_1099_),
    .C(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__nand3_1 _4655_ (.A(_1082_),
    .B(_1099_),
    .C(_1100_),
    .Y(_1102_));
 sky130_fd_sc_hd__a21oi_2 _4656_ (.A1(_1099_),
    .A2(_1100_),
    .B1(_1082_),
    .Y(_1103_));
 sky130_fd_sc_hd__a211oi_4 _4657_ (.A1(_1032_),
    .A2(_1035_),
    .B1(_1101_),
    .C1(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__o211a_1 _4658_ (.A1(_1101_),
    .A2(_1103_),
    .B1(_1032_),
    .C1(_1035_),
    .X(_1105_));
 sky130_fd_sc_hd__nor3_1 _4659_ (.A(_1071_),
    .B(_1104_),
    .C(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__or3_1 _4660_ (.A(_1071_),
    .B(_1104_),
    .C(_1105_),
    .X(_1107_));
 sky130_fd_sc_hd__o21ai_1 _4661_ (.A1(_1104_),
    .A2(_1105_),
    .B1(_1071_),
    .Y(_1108_));
 sky130_fd_sc_hd__o211a_1 _4662_ (.A1(_1037_),
    .A2(_1039_),
    .B1(_1107_),
    .C1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__a211oi_2 _4663_ (.A1(_1107_),
    .A2(_1108_),
    .B1(_1037_),
    .C1(_1039_),
    .Y(_1110_));
 sky130_fd_sc_hd__nor3_1 _4664_ (.A(_1002_),
    .B(_1109_),
    .C(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__or3_1 _4665_ (.A(_1002_),
    .B(_1109_),
    .C(_1110_),
    .X(_1112_));
 sky130_fd_sc_hd__o21ai_1 _4666_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1002_),
    .Y(_1113_));
 sky130_fd_sc_hd__o211a_1 _4667_ (.A1(_1041_),
    .A2(_1043_),
    .B1(_1112_),
    .C1(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__inv_2 _4668_ (.A(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__a211o_1 _4669_ (.A1(_1112_),
    .A2(_1113_),
    .B1(_1041_),
    .C1(_1043_),
    .X(_1116_));
 sky130_fd_sc_hd__nand2b_1 _4670_ (.A_N(_1114_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__a31o_1 _4671_ (.A1(_0925_),
    .A2(_0983_),
    .A3(_1047_),
    .B1(_1045_),
    .X(_1118_));
 sky130_fd_sc_hd__xor2_1 _4672_ (.A(_1117_),
    .B(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__or2_1 _4673_ (.A(_1051_),
    .B(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_1051_),
    .B(_1119_),
    .Y(_1121_));
 sky130_fd_sc_hd__and2_1 _4675_ (.A(_1120_),
    .B(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__a32o_1 _4676_ (.A1(_0933_),
    .A2(_0989_),
    .A3(_0990_),
    .B1(_1051_),
    .B2(_1052_),
    .X(_1123_));
 sky130_fd_sc_hd__a32o_1 _4677_ (.A1(_0993_),
    .A2(_1051_),
    .A3(_1052_),
    .B1(_1123_),
    .B2(_0987_),
    .X(_1124_));
 sky130_fd_sc_hd__or2_1 _4678_ (.A(_1122_),
    .B(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nand2_1 _4679_ (.A(_1122_),
    .B(_1124_),
    .Y(_1126_));
 sky130_fd_sc_hd__and3_1 _4680_ (.A(net208),
    .B(_1125_),
    .C(_1126_),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _4681_ (.A(_1048_),
    .B(_1117_),
    .X(_1127_));
 sky130_fd_sc_hd__a21oi_1 _4682_ (.A1(_0999_),
    .A2(_1070_),
    .B1(_1069_),
    .Y(_1128_));
 sky130_fd_sc_hd__a22oi_1 _4683_ (.A1(net141),
    .A2(net154),
    .B1(net151),
    .B2(net144),
    .Y(_1129_));
 sky130_fd_sc_hd__and4_1 _4684_ (.A(net141),
    .B(\ann.in_ff[2][0] ),
    .C(net154),
    .D(net151),
    .X(_1130_));
 sky130_fd_sc_hd__nor2_1 _4685_ (.A(_1129_),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__or2_1 _4686_ (.A(_1060_),
    .B(_1061_),
    .X(_1132_));
 sky130_fd_sc_hd__a22oi_1 _4687_ (.A1(net133),
    .A2(net161),
    .B1(net158),
    .B2(net136),
    .Y(_1133_));
 sky130_fd_sc_hd__and4_1 _4688_ (.A(net133),
    .B(net136),
    .C(net161),
    .D(net158),
    .X(_1134_));
 sky130_fd_sc_hd__and4bb_1 _4689_ (.A_N(_1133_),
    .B_N(_1134_),
    .C(net139),
    .D(net156),
    .X(_1135_));
 sky130_fd_sc_hd__o2bb2a_1 _4690_ (.A1_N(net139),
    .A2_N(net157),
    .B1(_1133_),
    .B2(_1134_),
    .X(_1136_));
 sky130_fd_sc_hd__nor2_1 _4691_ (.A(_1135_),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__and2_1 _4692_ (.A(_1132_),
    .B(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__xor2_1 _4693_ (.A(_1132_),
    .B(_1137_),
    .X(_1139_));
 sky130_fd_sc_hd__and2_1 _4694_ (.A(_1131_),
    .B(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__xnor2_1 _4695_ (.A(_1131_),
    .B(_1139_),
    .Y(_1141_));
 sky130_fd_sc_hd__a21oi_2 _4696_ (.A1(_1079_),
    .A2(_1081_),
    .B1(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__and3_1 _4697_ (.A(_1079_),
    .B(_1081_),
    .C(_1141_),
    .X(_1143_));
 sky130_fd_sc_hd__a211oi_2 _4698_ (.A1(_1064_),
    .A2(_1066_),
    .B1(_1142_),
    .C1(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__o211a_1 _4699_ (.A1(_1142_),
    .A2(_1143_),
    .B1(_1064_),
    .C1(_1066_),
    .X(_1145_));
 sky130_fd_sc_hd__or2_1 _4700_ (.A(_1074_),
    .B(_1075_),
    .X(_1146_));
 sky130_fd_sc_hd__a22oi_1 _4701_ (.A1(net125),
    .A2(net168),
    .B1(net166),
    .B2(net128),
    .Y(_1147_));
 sky130_fd_sc_hd__and4_1 _4702_ (.A(\ann.in_ff[2][7] ),
    .B(net128),
    .C(net168),
    .D(net166),
    .X(_1148_));
 sky130_fd_sc_hd__and4bb_1 _4703_ (.A_N(_1147_),
    .B_N(_1148_),
    .C(net130),
    .D(net164),
    .X(_1149_));
 sky130_fd_sc_hd__o2bb2a_1 _4704_ (.A1_N(net130),
    .A2_N(net164),
    .B1(_1147_),
    .B2(_1148_),
    .X(_1150_));
 sky130_fd_sc_hd__nor2_1 _4705_ (.A(_1149_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__o21ba_1 _4706_ (.A1(_1084_),
    .A2(_1085_),
    .B1_N(_1086_),
    .X(_1152_));
 sky130_fd_sc_hd__or3_1 _4707_ (.A(_1149_),
    .B(_1150_),
    .C(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__xnor2_2 _4708_ (.A(_1151_),
    .B(_1152_),
    .Y(_1154_));
 sky130_fd_sc_hd__nand2_1 _4709_ (.A(_1146_),
    .B(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__xor2_2 _4710_ (.A(_1146_),
    .B(_1154_),
    .X(_1156_));
 sky130_fd_sc_hd__a21bo_1 _4711_ (.A1(_1088_),
    .A2(_1096_),
    .B1_N(_1095_),
    .X(_1157_));
 sky130_fd_sc_hd__nand2_1 _4712_ (.A(net124),
    .B(net172),
    .Y(_1158_));
 sky130_fd_sc_hd__a22oi_2 _4713_ (.A1(net117),
    .A2(net176),
    .B1(net173),
    .B2(net121),
    .Y(_1159_));
 sky130_fd_sc_hd__and4_1 _4714_ (.A(net118),
    .B(net121),
    .C(net176),
    .D(net173),
    .X(_1160_));
 sky130_fd_sc_hd__nor2_1 _4715_ (.A(_1159_),
    .B(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__xnor2_2 _4716_ (.A(_1158_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__a21bo_1 _4717_ (.A1(_1090_),
    .A2(_1091_),
    .B1_N(_1092_),
    .X(_1163_));
 sky130_fd_sc_hd__and2_1 _4718_ (.A(net114),
    .B(net177),
    .X(_1164_));
 sky130_fd_sc_hd__a22o_1 _4719_ (.A1(net109),
    .A2(net181),
    .B1(net179),
    .B2(net111),
    .X(_1165_));
 sky130_fd_sc_hd__nand4_2 _4720_ (.A(net109),
    .B(net111),
    .C(net181),
    .D(net179),
    .Y(_1166_));
 sky130_fd_sc_hd__nand3_1 _4721_ (.A(_1164_),
    .B(_1165_),
    .C(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__a21o_1 _4722_ (.A1(_1165_),
    .A2(_1166_),
    .B1(_1164_),
    .X(_1168_));
 sky130_fd_sc_hd__nand3_2 _4723_ (.A(_1163_),
    .B(_1167_),
    .C(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__a21o_1 _4724_ (.A1(_1167_),
    .A2(_1168_),
    .B1(_1163_),
    .X(_1170_));
 sky130_fd_sc_hd__nand3_2 _4725_ (.A(_1162_),
    .B(_1169_),
    .C(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__a21o_1 _4726_ (.A1(_1169_),
    .A2(_1170_),
    .B1(_1162_),
    .X(_1172_));
 sky130_fd_sc_hd__nand3_4 _4727_ (.A(_1157_),
    .B(_1171_),
    .C(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__a21o_1 _4728_ (.A1(_1171_),
    .A2(_1172_),
    .B1(_1157_),
    .X(_1174_));
 sky130_fd_sc_hd__and3_1 _4729_ (.A(_1156_),
    .B(_1173_),
    .C(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__nand3_2 _4730_ (.A(_1156_),
    .B(_1173_),
    .C(_1174_),
    .Y(_1176_));
 sky130_fd_sc_hd__a21oi_1 _4731_ (.A1(_1173_),
    .A2(_1174_),
    .B1(_1156_),
    .Y(_1177_));
 sky130_fd_sc_hd__a211o_1 _4732_ (.A1(_1099_),
    .A2(_1102_),
    .B1(_1175_),
    .C1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__o211ai_2 _4733_ (.A1(_1175_),
    .A2(_1177_),
    .B1(_1099_),
    .C1(_1102_),
    .Y(_1179_));
 sky130_fd_sc_hd__or4bb_2 _4734_ (.A(_1144_),
    .B(_1145_),
    .C_N(_1178_),
    .D_N(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__a2bb2o_1 _4735_ (.A1_N(_1144_),
    .A2_N(_1145_),
    .B1(_1178_),
    .B2(_1179_),
    .X(_1181_));
 sky130_fd_sc_hd__o211a_1 _4736_ (.A1(_1104_),
    .A2(_1106_),
    .B1(_1180_),
    .C1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__a211oi_2 _4737_ (.A1(_1180_),
    .A2(_1181_),
    .B1(_1104_),
    .C1(_1106_),
    .Y(_1183_));
 sky130_fd_sc_hd__nor3_1 _4738_ (.A(_1128_),
    .B(_1182_),
    .C(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__or3_1 _4739_ (.A(_1128_),
    .B(_1182_),
    .C(_1183_),
    .X(_1185_));
 sky130_fd_sc_hd__o21ai_1 _4740_ (.A1(_1182_),
    .A2(_1183_),
    .B1(_1128_),
    .Y(_1186_));
 sky130_fd_sc_hd__o211a_1 _4741_ (.A1(_1109_),
    .A2(_1111_),
    .B1(_1185_),
    .C1(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__a211o_1 _4742_ (.A1(_1185_),
    .A2(_1186_),
    .B1(_1109_),
    .C1(_1111_),
    .X(_1188_));
 sky130_fd_sc_hd__nand2b_1 _4743_ (.A_N(_1187_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__a21oi_1 _4744_ (.A1(_1045_),
    .A2(_1116_),
    .B1(_1114_),
    .Y(_1190_));
 sky130_fd_sc_hd__xnor2_1 _4745_ (.A(_1189_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__nor2_1 _4746_ (.A(_1127_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__or2_1 _4747_ (.A(_1127_),
    .B(_1191_),
    .X(_1193_));
 sky130_fd_sc_hd__and2_1 _4748_ (.A(_1127_),
    .B(_1191_),
    .X(_1194_));
 sky130_fd_sc_hd__nor2_1 _4749_ (.A(_1192_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand2_1 _4750_ (.A(_1120_),
    .B(_1126_),
    .Y(_1196_));
 sky130_fd_sc_hd__xnor2_1 _4751_ (.A(_1195_),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__nor2_1 _4752_ (.A(net195),
    .B(_1197_),
    .Y(_0004_));
 sky130_fd_sc_hd__and3_1 _4753_ (.A(_1122_),
    .B(_1124_),
    .C(_1195_),
    .X(_1198_));
 sky130_fd_sc_hd__a21oi_1 _4754_ (.A1(_1120_),
    .A2(_1193_),
    .B1(_1194_),
    .Y(_1199_));
 sky130_fd_sc_hd__or3_1 _4755_ (.A(_1046_),
    .B(_1117_),
    .C(_1189_),
    .X(_1200_));
 sky130_fd_sc_hd__o21ai_1 _4756_ (.A1(_1142_),
    .A2(_1144_),
    .B1(_1130_),
    .Y(_1201_));
 sky130_fd_sc_hd__or3_1 _4757_ (.A(_1130_),
    .B(_1142_),
    .C(_1144_),
    .X(_1202_));
 sky130_fd_sc_hd__and2_1 _4758_ (.A(_1201_),
    .B(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(net144),
    .B(net149),
    .Y(_1204_));
 sky130_fd_sc_hd__a22oi_2 _4760_ (.A1(net138),
    .A2(net154),
    .B1(net152),
    .B2(net142),
    .Y(_1205_));
 sky130_fd_sc_hd__and4_1 _4761_ (.A(net138),
    .B(net142),
    .C(net154),
    .D(net152),
    .X(_1206_));
 sky130_fd_sc_hd__nor2_1 _4762_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__xnor2_1 _4763_ (.A(_1204_),
    .B(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__or2_1 _4764_ (.A(_1134_),
    .B(_1135_),
    .X(_1209_));
 sky130_fd_sc_hd__a22oi_1 _4765_ (.A1(net129),
    .A2(net161),
    .B1(net158),
    .B2(net132),
    .Y(_1210_));
 sky130_fd_sc_hd__and4_1 _4766_ (.A(net129),
    .B(net132),
    .C(net161),
    .D(net158),
    .X(_1211_));
 sky130_fd_sc_hd__and4bb_1 _4767_ (.A_N(_1210_),
    .B_N(_1211_),
    .C(net135),
    .D(net156),
    .X(_1212_));
 sky130_fd_sc_hd__o2bb2a_1 _4768_ (.A1_N(net135),
    .A2_N(net156),
    .B1(_1210_),
    .B2(_1211_),
    .X(_1213_));
 sky130_fd_sc_hd__nor2_1 _4769_ (.A(_1212_),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__and2_1 _4770_ (.A(_1209_),
    .B(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__xor2_1 _4771_ (.A(_1209_),
    .B(_1214_),
    .X(_1216_));
 sky130_fd_sc_hd__and2_1 _4772_ (.A(_1208_),
    .B(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__xnor2_1 _4773_ (.A(_1208_),
    .B(_1216_),
    .Y(_1218_));
 sky130_fd_sc_hd__a21o_2 _4774_ (.A1(_1153_),
    .A2(_1155_),
    .B1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__nand3_2 _4775_ (.A(_1153_),
    .B(_1155_),
    .C(_1218_),
    .Y(_1220_));
 sky130_fd_sc_hd__o211ai_4 _4776_ (.A1(_1138_),
    .A2(_1140_),
    .B1(_1219_),
    .C1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__a211o_1 _4777_ (.A1(_1219_),
    .A2(_1220_),
    .B1(_1138_),
    .C1(_1140_),
    .X(_1222_));
 sky130_fd_sc_hd__or2_1 _4778_ (.A(_1148_),
    .B(_1149_),
    .X(_1223_));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(net127),
    .B(net164),
    .Y(_1224_));
 sky130_fd_sc_hd__a22o_1 _4780_ (.A1(net123),
    .A2(net168),
    .B1(net166),
    .B2(net125),
    .X(_1225_));
 sky130_fd_sc_hd__and3_1 _4781_ (.A(net123),
    .B(net125),
    .C(net166),
    .X(_1226_));
 sky130_fd_sc_hd__a21bo_1 _4782_ (.A1(net168),
    .A2(_1226_),
    .B1_N(_1225_),
    .X(_1227_));
 sky130_fd_sc_hd__xor2_2 _4783_ (.A(_1224_),
    .B(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__o21ba_1 _4784_ (.A1(_1158_),
    .A2(_1159_),
    .B1_N(_1160_),
    .X(_1229_));
 sky130_fd_sc_hd__nand2b_1 _4785_ (.A_N(_1229_),
    .B(_1228_),
    .Y(_1230_));
 sky130_fd_sc_hd__xnor2_2 _4786_ (.A(_1228_),
    .B(_1229_),
    .Y(_1231_));
 sky130_fd_sc_hd__nand2_1 _4787_ (.A(_1223_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__xor2_2 _4788_ (.A(_1223_),
    .B(_1231_),
    .X(_1233_));
 sky130_fd_sc_hd__a21bo_1 _4789_ (.A1(_1162_),
    .A2(_1170_),
    .B1_N(_1169_),
    .X(_1234_));
 sky130_fd_sc_hd__a22oi_1 _4790_ (.A1(net114),
    .A2(net176),
    .B1(net173),
    .B2(net117),
    .Y(_1235_));
 sky130_fd_sc_hd__and4_1 _4791_ (.A(net115),
    .B(net117),
    .C(net176),
    .D(net173),
    .X(_1236_));
 sky130_fd_sc_hd__and4bb_1 _4792_ (.A_N(_1235_),
    .B_N(_1236_),
    .C(net120),
    .D(net172),
    .X(_1237_));
 sky130_fd_sc_hd__o2bb2a_1 _4793_ (.A1_N(net120),
    .A2_N(net172),
    .B1(_1235_),
    .B2(_1236_),
    .X(_1238_));
 sky130_fd_sc_hd__nor2_1 _4794_ (.A(_1237_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__a21bo_1 _4795_ (.A1(_1164_),
    .A2(_1165_),
    .B1_N(_1166_),
    .X(_1240_));
 sky130_fd_sc_hd__and2_1 _4796_ (.A(net111),
    .B(\ann.weight[2] ),
    .X(_1241_));
 sky130_fd_sc_hd__a22o_1 _4797_ (.A1(net107),
    .A2(net181),
    .B1(net179),
    .B2(net109),
    .X(_1242_));
 sky130_fd_sc_hd__nand4_1 _4798_ (.A(net107),
    .B(net109),
    .C(net181),
    .D(net179),
    .Y(_1243_));
 sky130_fd_sc_hd__nand3_1 _4799_ (.A(_1241_),
    .B(_1242_),
    .C(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__a21o_1 _4800_ (.A1(_1242_),
    .A2(_1243_),
    .B1(_1241_),
    .X(_1245_));
 sky130_fd_sc_hd__nand3_1 _4801_ (.A(_1240_),
    .B(_1244_),
    .C(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a21o_1 _4802_ (.A1(_1244_),
    .A2(_1245_),
    .B1(_1240_),
    .X(_1247_));
 sky130_fd_sc_hd__nand3_2 _4803_ (.A(_1239_),
    .B(_1246_),
    .C(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__a21o_1 _4804_ (.A1(_1246_),
    .A2(_1247_),
    .B1(_1239_),
    .X(_1249_));
 sky130_fd_sc_hd__nand3_4 _4805_ (.A(_1234_),
    .B(_1248_),
    .C(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__a21o_1 _4806_ (.A1(_1248_),
    .A2(_1249_),
    .B1(_1234_),
    .X(_1251_));
 sky130_fd_sc_hd__and3_1 _4807_ (.A(_1233_),
    .B(_1250_),
    .C(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__nand3_2 _4808_ (.A(_1233_),
    .B(_1250_),
    .C(_1251_),
    .Y(_1253_));
 sky130_fd_sc_hd__a21oi_2 _4809_ (.A1(_1250_),
    .A2(_1251_),
    .B1(_1233_),
    .Y(_1254_));
 sky130_fd_sc_hd__a211oi_2 _4810_ (.A1(_1173_),
    .A2(_1176_),
    .B1(_1252_),
    .C1(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__a211o_1 _4811_ (.A1(_1173_),
    .A2(_1176_),
    .B1(_1252_),
    .C1(_1254_),
    .X(_1256_));
 sky130_fd_sc_hd__o211ai_2 _4812_ (.A1(_1252_),
    .A2(_1254_),
    .B1(_1173_),
    .C1(_1176_),
    .Y(_1257_));
 sky130_fd_sc_hd__and4_2 _4813_ (.A(_1221_),
    .B(_1222_),
    .C(_1256_),
    .D(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__a22oi_2 _4814_ (.A1(_1221_),
    .A2(_1222_),
    .B1(_1256_),
    .B2(_1257_),
    .Y(_1259_));
 sky130_fd_sc_hd__a211o_2 _4815_ (.A1(_1178_),
    .A2(_1180_),
    .B1(_1258_),
    .C1(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__o211ai_2 _4816_ (.A1(_1258_),
    .A2(_1259_),
    .B1(_1178_),
    .C1(_1180_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand3_2 _4817_ (.A(_1203_),
    .B(_1260_),
    .C(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__a21o_1 _4818_ (.A1(_1260_),
    .A2(_1261_),
    .B1(_1203_),
    .X(_1263_));
 sky130_fd_sc_hd__o211a_1 _4819_ (.A1(_1182_),
    .A2(_1184_),
    .B1(_1262_),
    .C1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__a211o_1 _4820_ (.A1(_1262_),
    .A2(_1263_),
    .B1(_1182_),
    .C1(_1184_),
    .X(_1265_));
 sky130_fd_sc_hd__and2b_1 _4821_ (.A_N(_1264_),
    .B(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__a21o_1 _4822_ (.A1(_1114_),
    .A2(_1188_),
    .B1(_1187_),
    .X(_1267_));
 sky130_fd_sc_hd__xnor2_2 _4823_ (.A(_1266_),
    .B(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__nor2_1 _4824_ (.A(_1200_),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__or2_1 _4825_ (.A(_1200_),
    .B(_1268_),
    .X(_1270_));
 sky130_fd_sc_hd__xor2_1 _4826_ (.A(_1200_),
    .B(_1268_),
    .X(_1271_));
 sky130_fd_sc_hd__or3_1 _4827_ (.A(_1198_),
    .B(_1199_),
    .C(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__o21ai_1 _4828_ (.A1(_1198_),
    .A2(_1199_),
    .B1(_1271_),
    .Y(_1273_));
 sky130_fd_sc_hd__and3_1 _4829_ (.A(net208),
    .B(_1272_),
    .C(_1273_),
    .X(_0005_));
 sky130_fd_sc_hd__nand2_1 _4830_ (.A(_1270_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__or3b_1 _4831_ (.A(_1115_),
    .B(_1189_),
    .C_N(_1266_),
    .X(_1275_));
 sky130_fd_sc_hd__nand2_8 _4832_ (.A(net144),
    .B(net147),
    .Y(_1276_));
 sky130_fd_sc_hd__o21ba_1 _4833_ (.A1(_1204_),
    .A2(_1205_),
    .B1_N(_1206_),
    .X(_1277_));
 sky130_fd_sc_hd__nor2_1 _4834_ (.A(_1276_),
    .B(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__xnor2_1 _4835_ (.A(_1276_),
    .B(_1277_),
    .Y(_1279_));
 sky130_fd_sc_hd__a21oi_1 _4836_ (.A1(_1219_),
    .A2(_1221_),
    .B1(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__and3_1 _4837_ (.A(_1219_),
    .B(_1221_),
    .C(_1279_),
    .X(_1281_));
 sky130_fd_sc_hd__or2_1 _4838_ (.A(_1280_),
    .B(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__a22oi_1 _4839_ (.A1(net135),
    .A2(net153),
    .B1(net151),
    .B2(net138),
    .Y(_1283_));
 sky130_fd_sc_hd__and4_1 _4840_ (.A(net135),
    .B(net138),
    .C(net154),
    .D(net151),
    .X(_1284_));
 sky130_fd_sc_hd__nor2_1 _4841_ (.A(_1283_),
    .B(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__a21oi_1 _4842_ (.A1(net142),
    .A2(net149),
    .B1(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__and3_1 _4843_ (.A(net142),
    .B(net149),
    .C(_1285_),
    .X(_1287_));
 sky130_fd_sc_hd__nor2_1 _4844_ (.A(_1286_),
    .B(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__or2_1 _4845_ (.A(_1211_),
    .B(_1212_),
    .X(_1289_));
 sky130_fd_sc_hd__nand2_1 _4846_ (.A(net132),
    .B(net156),
    .Y(_1290_));
 sky130_fd_sc_hd__a22o_1 _4847_ (.A1(net127),
    .A2(net161),
    .B1(net158),
    .B2(net129),
    .X(_1291_));
 sky130_fd_sc_hd__and3_1 _4848_ (.A(net127),
    .B(net129),
    .C(net158),
    .X(_1292_));
 sky130_fd_sc_hd__a21bo_1 _4849_ (.A1(net161),
    .A2(_1292_),
    .B1_N(_1291_),
    .X(_1293_));
 sky130_fd_sc_hd__xor2_1 _4850_ (.A(_1290_),
    .B(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__and2_1 _4851_ (.A(_1289_),
    .B(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__xor2_1 _4852_ (.A(_1289_),
    .B(_1294_),
    .X(_1296_));
 sky130_fd_sc_hd__xnor2_1 _4853_ (.A(_1288_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__a21o_2 _4854_ (.A1(_1230_),
    .A2(_1232_),
    .B1(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__nand3_2 _4855_ (.A(_1230_),
    .B(_1232_),
    .C(_1297_),
    .Y(_1299_));
 sky130_fd_sc_hd__o211ai_4 _4856_ (.A1(_1215_),
    .A2(_1217_),
    .B1(_1298_),
    .C1(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__a211o_1 _4857_ (.A1(_1298_),
    .A2(_1299_),
    .B1(_1215_),
    .C1(_1217_),
    .X(_1301_));
 sky130_fd_sc_hd__a32o_1 _4858_ (.A1(net127),
    .A2(net164),
    .A3(_1225_),
    .B1(_1226_),
    .B2(net168),
    .X(_1302_));
 sky130_fd_sc_hd__a22o_1 _4859_ (.A1(net120),
    .A2(net168),
    .B1(net166),
    .B2(net123),
    .X(_1303_));
 sky130_fd_sc_hd__nand4_2 _4860_ (.A(net120),
    .B(net123),
    .C(net168),
    .D(net166),
    .Y(_1304_));
 sky130_fd_sc_hd__nand4_2 _4861_ (.A(net125),
    .B(net164),
    .C(_1303_),
    .D(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__a22o_1 _4862_ (.A1(net125),
    .A2(net164),
    .B1(_1303_),
    .B2(_1304_),
    .X(_1306_));
 sky130_fd_sc_hd__o211a_1 _4863_ (.A1(_1236_),
    .A2(_1237_),
    .B1(_1305_),
    .C1(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__a211o_1 _4864_ (.A1(_1305_),
    .A2(_1306_),
    .B1(_1236_),
    .C1(_1237_),
    .X(_1308_));
 sky130_fd_sc_hd__nand2b_1 _4865_ (.A_N(_1307_),
    .B(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__xnor2_1 _4866_ (.A(_1302_),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__a21bo_1 _4867_ (.A1(_1239_),
    .A2(_1247_),
    .B1_N(_1246_),
    .X(_1311_));
 sky130_fd_sc_hd__a22oi_1 _4868_ (.A1(net112),
    .A2(net176),
    .B1(net173),
    .B2(net114),
    .Y(_1312_));
 sky130_fd_sc_hd__and4_1 _4869_ (.A(net112),
    .B(net115),
    .C(net176),
    .D(net173),
    .X(_1313_));
 sky130_fd_sc_hd__and4bb_1 _4870_ (.A_N(_1312_),
    .B_N(_1313_),
    .C(net117),
    .D(net172),
    .X(_1314_));
 sky130_fd_sc_hd__o2bb2a_1 _4871_ (.A1_N(net117),
    .A2_N(net172),
    .B1(_1312_),
    .B2(_1313_),
    .X(_1315_));
 sky130_fd_sc_hd__nor2_1 _4872_ (.A(_1314_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__a21bo_1 _4873_ (.A1(_1241_),
    .A2(_1242_),
    .B1_N(_1243_),
    .X(_1317_));
 sky130_fd_sc_hd__and2_1 _4874_ (.A(net109),
    .B(\ann.weight[2] ),
    .X(_1318_));
 sky130_fd_sc_hd__a22o_1 _4875_ (.A1(net105),
    .A2(net181),
    .B1(net179),
    .B2(net107),
    .X(_1319_));
 sky130_fd_sc_hd__nand4_2 _4876_ (.A(net105),
    .B(net107),
    .C(net181),
    .D(net179),
    .Y(_1320_));
 sky130_fd_sc_hd__nand3_1 _4877_ (.A(_1318_),
    .B(_1319_),
    .C(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__a21o_1 _4878_ (.A1(_1319_),
    .A2(_1320_),
    .B1(_1318_),
    .X(_1322_));
 sky130_fd_sc_hd__nand3_1 _4879_ (.A(_1317_),
    .B(_1321_),
    .C(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__a21o_1 _4880_ (.A1(_1321_),
    .A2(_1322_),
    .B1(_1317_),
    .X(_1324_));
 sky130_fd_sc_hd__nand3_1 _4881_ (.A(_1316_),
    .B(_1323_),
    .C(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__a21o_1 _4882_ (.A1(_1323_),
    .A2(_1324_),
    .B1(_1316_),
    .X(_1326_));
 sky130_fd_sc_hd__nand3_2 _4883_ (.A(_1311_),
    .B(_1325_),
    .C(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__a21o_1 _4884_ (.A1(_1325_),
    .A2(_1326_),
    .B1(_1311_),
    .X(_1328_));
 sky130_fd_sc_hd__and3_1 _4885_ (.A(_1310_),
    .B(_1327_),
    .C(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__nand3_1 _4886_ (.A(_1310_),
    .B(_1327_),
    .C(_1328_),
    .Y(_1330_));
 sky130_fd_sc_hd__a21oi_2 _4887_ (.A1(_1327_),
    .A2(_1328_),
    .B1(_1310_),
    .Y(_1331_));
 sky130_fd_sc_hd__a211o_2 _4888_ (.A1(_1250_),
    .A2(_1253_),
    .B1(_1329_),
    .C1(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__inv_2 _4889_ (.A(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__o211ai_4 _4890_ (.A1(_1329_),
    .A2(_1331_),
    .B1(_1250_),
    .C1(_1253_),
    .Y(_1334_));
 sky130_fd_sc_hd__and4_1 _4891_ (.A(_1300_),
    .B(_1301_),
    .C(_1332_),
    .D(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__nand4_1 _4892_ (.A(_1300_),
    .B(_1301_),
    .C(_1332_),
    .D(_1334_),
    .Y(_1336_));
 sky130_fd_sc_hd__a22o_1 _4893_ (.A1(_1300_),
    .A2(_1301_),
    .B1(_1332_),
    .B2(_1334_),
    .X(_1337_));
 sky130_fd_sc_hd__o211a_1 _4894_ (.A1(_1255_),
    .A2(_1258_),
    .B1(_1336_),
    .C1(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__a211oi_2 _4895_ (.A1(_1336_),
    .A2(_1337_),
    .B1(_1255_),
    .C1(_1258_),
    .Y(_1339_));
 sky130_fd_sc_hd__nor3_2 _4896_ (.A(_1282_),
    .B(_1338_),
    .C(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__o21a_1 _4897_ (.A1(_1338_),
    .A2(_1339_),
    .B1(_1282_),
    .X(_1341_));
 sky130_fd_sc_hd__a211oi_1 _4898_ (.A1(_1260_),
    .A2(_1262_),
    .B1(_1340_),
    .C1(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__a211o_1 _4899_ (.A1(_1260_),
    .A2(_1262_),
    .B1(_1340_),
    .C1(_1341_),
    .X(_1343_));
 sky130_fd_sc_hd__o211a_1 _4900_ (.A1(_1340_),
    .A2(_1341_),
    .B1(_1260_),
    .C1(_1262_),
    .X(_1344_));
 sky130_fd_sc_hd__or3_4 _4901_ (.A(_1201_),
    .B(_1342_),
    .C(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__o21ai_1 _4902_ (.A1(_1342_),
    .A2(_1344_),
    .B1(_1201_),
    .Y(_1346_));
 sky130_fd_sc_hd__and2_1 _4903_ (.A(_1345_),
    .B(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a21oi_1 _4904_ (.A1(_1187_),
    .A2(_1265_),
    .B1(_1264_),
    .Y(_1348_));
 sky130_fd_sc_hd__nand3_1 _4905_ (.A(_1345_),
    .B(_1346_),
    .C(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__a21o_1 _4906_ (.A1(_1345_),
    .A2(_1346_),
    .B1(_1348_),
    .X(_1350_));
 sky130_fd_sc_hd__a21oi_1 _4907_ (.A1(_1349_),
    .A2(_1350_),
    .B1(_1275_),
    .Y(_1351_));
 sky130_fd_sc_hd__nand3_2 _4908_ (.A(_1275_),
    .B(_1349_),
    .C(_1350_),
    .Y(_1352_));
 sky130_fd_sc_hd__nand2b_1 _4909_ (.A_N(_1351_),
    .B(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__and3_1 _4910_ (.A(_1270_),
    .B(_1273_),
    .C(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__a211oi_2 _4911_ (.A1(_1274_),
    .A2(_1352_),
    .B1(_1354_),
    .C1(net195),
    .Y(_0006_));
 sky130_fd_sc_hd__a21o_1 _4912_ (.A1(_1269_),
    .A2(_1352_),
    .B1(_1351_),
    .X(_1355_));
 sky130_fd_sc_hd__and3b_1 _4913_ (.A_N(_1351_),
    .B(_1352_),
    .C(_1271_),
    .X(_1356_));
 sky130_fd_sc_hd__and2_1 _4914_ (.A(_1199_),
    .B(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__and4_1 _4915_ (.A(_1122_),
    .B(_1124_),
    .C(_1195_),
    .D(_1356_),
    .X(_1358_));
 sky130_fd_sc_hd__nand2_4 _4916_ (.A(net142),
    .B(net146),
    .Y(_1359_));
 sky130_fd_sc_hd__nor2_8 _4917_ (.A(_1276_),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__or2_1 _4918_ (.A(_1276_),
    .B(_1359_),
    .X(_1361_));
 sky130_fd_sc_hd__and2_2 _4919_ (.A(_1276_),
    .B(_1359_),
    .X(_1362_));
 sky130_fd_sc_hd__nor2_8 _4920_ (.A(_1360_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__o21a_1 _4921_ (.A1(_1284_),
    .A2(_1287_),
    .B1(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__nor3_1 _4922_ (.A(_1284_),
    .B(_1287_),
    .C(_1363_),
    .Y(_1365_));
 sky130_fd_sc_hd__nor2_1 _4923_ (.A(_1364_),
    .B(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__nand2_2 _4924_ (.A(_1278_),
    .B(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__or2_1 _4925_ (.A(_1278_),
    .B(_1366_),
    .X(_1368_));
 sky130_fd_sc_hd__nand2_1 _4926_ (.A(_1367_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__nand2_1 _4927_ (.A(_1298_),
    .B(_1300_),
    .Y(_1370_));
 sky130_fd_sc_hd__a21oi_2 _4928_ (.A1(_1298_),
    .A2(_1300_),
    .B1(_1369_),
    .Y(_1371_));
 sky130_fd_sc_hd__xor2_1 _4929_ (.A(_1369_),
    .B(_1370_),
    .X(_1372_));
 sky130_fd_sc_hd__a21oi_1 _4930_ (.A1(_1288_),
    .A2(_1296_),
    .B1(_1295_),
    .Y(_1373_));
 sky130_fd_sc_hd__a22oi_1 _4931_ (.A1(net132),
    .A2(net154),
    .B1(net152),
    .B2(net135),
    .Y(_1374_));
 sky130_fd_sc_hd__and4_1 _4932_ (.A(net132),
    .B(net135),
    .C(net154),
    .D(net152),
    .X(_1375_));
 sky130_fd_sc_hd__nor2_1 _4933_ (.A(_1374_),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_1 _4934_ (.A(net138),
    .B(net149),
    .Y(_1377_));
 sky130_fd_sc_hd__and3_1 _4935_ (.A(net138),
    .B(net149),
    .C(_1376_),
    .X(_1378_));
 sky130_fd_sc_hd__xnor2_1 _4936_ (.A(_1376_),
    .B(_1377_),
    .Y(_1379_));
 sky130_fd_sc_hd__a32o_1 _4937_ (.A1(net132),
    .A2(net156),
    .A3(_1291_),
    .B1(_1292_),
    .B2(net161),
    .X(_1380_));
 sky130_fd_sc_hd__and2_1 _4938_ (.A(net129),
    .B(net156),
    .X(_1381_));
 sky130_fd_sc_hd__a22o_1 _4939_ (.A1(net125),
    .A2(net161),
    .B1(net158),
    .B2(net127),
    .X(_1382_));
 sky130_fd_sc_hd__nand4_1 _4940_ (.A(net125),
    .B(net127),
    .C(net161),
    .D(net158),
    .Y(_1383_));
 sky130_fd_sc_hd__nand3_1 _4941_ (.A(_1381_),
    .B(_1382_),
    .C(_1383_),
    .Y(_1384_));
 sky130_fd_sc_hd__a21o_1 _4942_ (.A1(_1382_),
    .A2(_1383_),
    .B1(_1381_),
    .X(_1385_));
 sky130_fd_sc_hd__nand3_2 _4943_ (.A(_1380_),
    .B(_1384_),
    .C(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__a21o_1 _4944_ (.A1(_1384_),
    .A2(_1385_),
    .B1(_1380_),
    .X(_1387_));
 sky130_fd_sc_hd__nand3_1 _4945_ (.A(_1379_),
    .B(_1386_),
    .C(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__a21o_1 _4946_ (.A1(_1386_),
    .A2(_1387_),
    .B1(_1379_),
    .X(_1389_));
 sky130_fd_sc_hd__a21o_1 _4947_ (.A1(_1302_),
    .A2(_1308_),
    .B1(_1307_),
    .X(_1390_));
 sky130_fd_sc_hd__and3_1 _4948_ (.A(_1388_),
    .B(_1389_),
    .C(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__a21oi_1 _4949_ (.A1(_1388_),
    .A2(_1389_),
    .B1(_1390_),
    .Y(_1392_));
 sky130_fd_sc_hd__nor2_1 _4950_ (.A(_1391_),
    .B(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__xnor2_1 _4951_ (.A(_1373_),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__nand2_1 _4952_ (.A(_1304_),
    .B(_1305_),
    .Y(_1395_));
 sky130_fd_sc_hd__a22o_1 _4953_ (.A1(net118),
    .A2(net168),
    .B1(net166),
    .B2(net121),
    .X(_1396_));
 sky130_fd_sc_hd__nand4_2 _4954_ (.A(net118),
    .B(net121),
    .C(net168),
    .D(net166),
    .Y(_1397_));
 sky130_fd_sc_hd__nand4_2 _4955_ (.A(net123),
    .B(net164),
    .C(_1396_),
    .D(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__a22o_1 _4956_ (.A1(net123),
    .A2(net164),
    .B1(_1396_),
    .B2(_1397_),
    .X(_1399_));
 sky130_fd_sc_hd__o211a_1 _4957_ (.A1(_1313_),
    .A2(_1314_),
    .B1(_1398_),
    .C1(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__a211o_1 _4958_ (.A1(_1398_),
    .A2(_1399_),
    .B1(_1313_),
    .C1(_1314_),
    .X(_1401_));
 sky130_fd_sc_hd__nand2b_1 _4959_ (.A_N(_1400_),
    .B(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__xnor2_2 _4960_ (.A(_1395_),
    .B(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__a21bo_1 _4961_ (.A1(_1316_),
    .A2(_1324_),
    .B1_N(_1323_),
    .X(_1404_));
 sky130_fd_sc_hd__a22oi_1 _4962_ (.A1(net110),
    .A2(net175),
    .B1(net174),
    .B2(net113),
    .Y(_1405_));
 sky130_fd_sc_hd__and4_1 _4963_ (.A(net110),
    .B(net113),
    .C(net175),
    .D(net174),
    .X(_1406_));
 sky130_fd_sc_hd__and4bb_1 _4964_ (.A_N(_1405_),
    .B_N(_1406_),
    .C(net116),
    .D(net171),
    .X(_1407_));
 sky130_fd_sc_hd__o2bb2a_1 _4965_ (.A1_N(net116),
    .A2_N(net171),
    .B1(_1405_),
    .B2(_1406_),
    .X(_1408_));
 sky130_fd_sc_hd__nor2_1 _4966_ (.A(_1407_),
    .B(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__a21bo_1 _4967_ (.A1(_1318_),
    .A2(_1319_),
    .B1_N(_1320_),
    .X(_1410_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(net108),
    .B(net177),
    .Y(_1411_));
 sky130_fd_sc_hd__o21ai_1 _4969_ (.A1(net180),
    .A2(net178),
    .B1(net106),
    .Y(_1412_));
 sky130_fd_sc_hd__o21a_1 _4970_ (.A1(net181),
    .A2(net178),
    .B1(net106),
    .X(_1413_));
 sky130_fd_sc_hd__and3_1 _4971_ (.A(net106),
    .B(net181),
    .C(net178),
    .X(_1414_));
 sky130_fd_sc_hd__o21ai_1 _4972_ (.A1(_1412_),
    .A2(_1414_),
    .B1(_1411_),
    .Y(_1415_));
 sky130_fd_sc_hd__or3_1 _4973_ (.A(_1411_),
    .B(_1412_),
    .C(_1414_),
    .X(_1416_));
 sky130_fd_sc_hd__nand3_1 _4974_ (.A(_1410_),
    .B(_1415_),
    .C(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__a21o_1 _4975_ (.A1(_1415_),
    .A2(_1416_),
    .B1(_1410_),
    .X(_1418_));
 sky130_fd_sc_hd__nand3_2 _4976_ (.A(_1409_),
    .B(_1417_),
    .C(_1418_),
    .Y(_1419_));
 sky130_fd_sc_hd__a21o_1 _4977_ (.A1(_1417_),
    .A2(_1418_),
    .B1(_1409_),
    .X(_1420_));
 sky130_fd_sc_hd__nand3_1 _4978_ (.A(_1404_),
    .B(_1419_),
    .C(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__a21o_1 _4979_ (.A1(_1419_),
    .A2(_1420_),
    .B1(_1404_),
    .X(_1422_));
 sky130_fd_sc_hd__and3_1 _4980_ (.A(_1403_),
    .B(_1421_),
    .C(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__a21oi_1 _4981_ (.A1(_1421_),
    .A2(_1422_),
    .B1(_1403_),
    .Y(_1424_));
 sky130_fd_sc_hd__a211o_1 _4982_ (.A1(_1327_),
    .A2(_1330_),
    .B1(_1423_),
    .C1(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__o211ai_2 _4983_ (.A1(_1423_),
    .A2(_1424_),
    .B1(_1327_),
    .C1(_1330_),
    .Y(_1426_));
 sky130_fd_sc_hd__nand3_1 _4984_ (.A(_1394_),
    .B(_1425_),
    .C(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__a21o_1 _4985_ (.A1(_1425_),
    .A2(_1426_),
    .B1(_1394_),
    .X(_1428_));
 sky130_fd_sc_hd__o211a_1 _4986_ (.A1(_1333_),
    .A2(_1335_),
    .B1(_1427_),
    .C1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__a211oi_2 _4987_ (.A1(_1427_),
    .A2(_1428_),
    .B1(_1333_),
    .C1(_1335_),
    .Y(_1430_));
 sky130_fd_sc_hd__or3_1 _4988_ (.A(_1372_),
    .B(_1429_),
    .C(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__o21ai_1 _4989_ (.A1(_1429_),
    .A2(_1430_),
    .B1(_1372_),
    .Y(_1432_));
 sky130_fd_sc_hd__o211a_1 _4990_ (.A1(_1338_),
    .A2(_1340_),
    .B1(_1431_),
    .C1(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__a211oi_2 _4991_ (.A1(_1431_),
    .A2(_1432_),
    .B1(_1338_),
    .C1(_1340_),
    .Y(_1434_));
 sky130_fd_sc_hd__nor3b_2 _4992_ (.A(_1433_),
    .B(_1434_),
    .C_N(_1280_),
    .Y(_1435_));
 sky130_fd_sc_hd__o21ba_1 _4993_ (.A1(_1433_),
    .A2(_1434_),
    .B1_N(_1280_),
    .X(_1436_));
 sky130_fd_sc_hd__a211oi_2 _4994_ (.A1(_1343_),
    .A2(_1345_),
    .B1(_1435_),
    .C1(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__a211o_1 _4995_ (.A1(_1343_),
    .A2(_1345_),
    .B1(_1435_),
    .C1(_1436_),
    .X(_1438_));
 sky130_fd_sc_hd__o211ai_2 _4996_ (.A1(_1435_),
    .A2(_1436_),
    .B1(_1343_),
    .C1(_1345_),
    .Y(_1439_));
 sky130_fd_sc_hd__and4_1 _4997_ (.A(_1264_),
    .B(_1347_),
    .C(_1438_),
    .D(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__nand4_1 _4998_ (.A(_1264_),
    .B(_1347_),
    .C(_1438_),
    .D(_1439_),
    .Y(_1441_));
 sky130_fd_sc_hd__a22oi_1 _4999_ (.A1(_1264_),
    .A2(_1347_),
    .B1(_1438_),
    .B2(_1439_),
    .Y(_1442_));
 sky130_fd_sc_hd__nor2_1 _5000_ (.A(_1440_),
    .B(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__and3_1 _5001_ (.A(_1187_),
    .B(_1266_),
    .C(_1347_),
    .X(_1444_));
 sky130_fd_sc_hd__nand3_1 _5002_ (.A(_1187_),
    .B(_1266_),
    .C(_1347_),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _5003_ (.A(_1443_),
    .B(_1444_),
    .Y(_1446_));
 sky130_fd_sc_hd__xnor2_1 _5004_ (.A(_1443_),
    .B(_1445_),
    .Y(_1447_));
 sky130_fd_sc_hd__or4_1 _5005_ (.A(_1355_),
    .B(_1357_),
    .C(_1358_),
    .D(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__o31ai_2 _5006_ (.A1(_1355_),
    .A2(_1357_),
    .A3(_1358_),
    .B1(_1447_),
    .Y(_1449_));
 sky130_fd_sc_hd__and3_1 _5007_ (.A(net208),
    .B(_1448_),
    .C(_1449_),
    .X(_0007_));
 sky130_fd_sc_hd__o21ba_1 _5008_ (.A1(_1372_),
    .A2(_1430_),
    .B1_N(_1429_),
    .X(_1450_));
 sky130_fd_sc_hd__o21bai_2 _5009_ (.A1(_1373_),
    .A2(_1392_),
    .B1_N(_1391_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_2 _5010_ (.A(net138),
    .B(net146),
    .Y(_1452_));
 sky130_fd_sc_hd__o21ai_4 _5011_ (.A1(net138),
    .A2(net142),
    .B1(net146),
    .Y(_1453_));
 sky130_fd_sc_hd__and3_1 _5012_ (.A(net138),
    .B(net142),
    .C(net146),
    .X(_1454_));
 sky130_fd_sc_hd__nor2_2 _5013_ (.A(_1453_),
    .B(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__xnor2_4 _5014_ (.A(_1276_),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__o21ai_1 _5015_ (.A1(_1375_),
    .A2(_1378_),
    .B1(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__inv_2 _5016_ (.A(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__nor3_1 _5017_ (.A(_1375_),
    .B(_1378_),
    .C(_1456_),
    .Y(_1459_));
 sky130_fd_sc_hd__nor2_1 _5018_ (.A(_1458_),
    .B(_1459_),
    .Y(_1460_));
 sky130_fd_sc_hd__nor2_1 _5019_ (.A(_1360_),
    .B(_1364_),
    .Y(_1461_));
 sky130_fd_sc_hd__xnor2_2 _5020_ (.A(_1460_),
    .B(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__xnor2_2 _5021_ (.A(_1451_),
    .B(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__nor2_1 _5022_ (.A(_1367_),
    .B(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__xor2_2 _5023_ (.A(_1367_),
    .B(_1463_),
    .X(_1465_));
 sky130_fd_sc_hd__a21bo_1 _5024_ (.A1(_1394_),
    .A2(_1426_),
    .B1_N(_1425_),
    .X(_1466_));
 sky130_fd_sc_hd__nand2_2 _5025_ (.A(_1386_),
    .B(_1388_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(net135),
    .B(net149),
    .Y(_1468_));
 sky130_fd_sc_hd__a22o_1 _5027_ (.A1(net129),
    .A2(net153),
    .B1(net151),
    .B2(net132),
    .X(_1469_));
 sky130_fd_sc_hd__and3_1 _5028_ (.A(net129),
    .B(net132),
    .C(net151),
    .X(_1470_));
 sky130_fd_sc_hd__a21bo_1 _5029_ (.A1(net153),
    .A2(_1470_),
    .B1_N(_1469_),
    .X(_1471_));
 sky130_fd_sc_hd__xor2_1 _5030_ (.A(_1468_),
    .B(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__a21bo_1 _5031_ (.A1(_1381_),
    .A2(_1382_),
    .B1_N(_1383_),
    .X(_1473_));
 sky130_fd_sc_hd__and2_1 _5032_ (.A(net127),
    .B(net157),
    .X(_1474_));
 sky130_fd_sc_hd__a22o_1 _5033_ (.A1(net124),
    .A2(net163),
    .B1(net160),
    .B2(net125),
    .X(_1475_));
 sky130_fd_sc_hd__nand4_1 _5034_ (.A(net124),
    .B(net125),
    .C(net163),
    .D(net160),
    .Y(_1476_));
 sky130_fd_sc_hd__nand3_1 _5035_ (.A(_1474_),
    .B(_1475_),
    .C(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__a21o_1 _5036_ (.A1(_1475_),
    .A2(_1476_),
    .B1(_1474_),
    .X(_1478_));
 sky130_fd_sc_hd__nand3_1 _5037_ (.A(_1473_),
    .B(_1477_),
    .C(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__a21o_1 _5038_ (.A1(_1477_),
    .A2(_1478_),
    .B1(_1473_),
    .X(_1480_));
 sky130_fd_sc_hd__nand3_1 _5039_ (.A(_1472_),
    .B(_1479_),
    .C(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__a21o_1 _5040_ (.A1(_1479_),
    .A2(_1480_),
    .B1(_1472_),
    .X(_1482_));
 sky130_fd_sc_hd__a21o_1 _5041_ (.A1(_1395_),
    .A2(_1401_),
    .B1(_1400_),
    .X(_1483_));
 sky130_fd_sc_hd__and3_1 _5042_ (.A(_1481_),
    .B(_1482_),
    .C(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__a21o_1 _5043_ (.A1(_1481_),
    .A2(_1482_),
    .B1(_1483_),
    .X(_1485_));
 sky130_fd_sc_hd__and2b_1 _5044_ (.A_N(_1484_),
    .B(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__xor2_2 _5045_ (.A(_1467_),
    .B(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__a21boi_2 _5046_ (.A1(_1403_),
    .A2(_1422_),
    .B1_N(_1421_),
    .Y(_1488_));
 sky130_fd_sc_hd__nand2_2 _5047_ (.A(_1397_),
    .B(_1398_),
    .Y(_1489_));
 sky130_fd_sc_hd__a22o_1 _5048_ (.A1(net116),
    .A2(net170),
    .B1(net167),
    .B2(net119),
    .X(_1490_));
 sky130_fd_sc_hd__nand4_2 _5049_ (.A(net116),
    .B(net119),
    .C(net170),
    .D(net167),
    .Y(_1491_));
 sky130_fd_sc_hd__nand4_2 _5050_ (.A(net122),
    .B(net165),
    .C(_1490_),
    .D(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__a22o_1 _5051_ (.A1(net122),
    .A2(net165),
    .B1(_1490_),
    .B2(_1491_),
    .X(_1493_));
 sky130_fd_sc_hd__o211a_1 _5052_ (.A1(_1406_),
    .A2(_1407_),
    .B1(_1492_),
    .C1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__a211o_1 _5053_ (.A1(_1492_),
    .A2(_1493_),
    .B1(_1406_),
    .C1(_1407_),
    .X(_1495_));
 sky130_fd_sc_hd__nand2b_1 _5054_ (.A_N(_1494_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__xnor2_2 _5055_ (.A(_1489_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__a21bo_1 _5056_ (.A1(_1409_),
    .A2(_1418_),
    .B1_N(_1417_),
    .X(_1498_));
 sky130_fd_sc_hd__nand2_1 _5057_ (.A(net113),
    .B(net171),
    .Y(_1499_));
 sky130_fd_sc_hd__a22o_1 _5058_ (.A1(net108),
    .A2(net175),
    .B1(net174),
    .B2(net110),
    .X(_1500_));
 sky130_fd_sc_hd__and3_1 _5059_ (.A(net108),
    .B(net110),
    .C(net174),
    .X(_1501_));
 sky130_fd_sc_hd__and4_1 _5060_ (.A(net108),
    .B(net110),
    .C(net175),
    .D(net174),
    .X(_1502_));
 sky130_fd_sc_hd__a21bo_1 _5061_ (.A1(net175),
    .A2(_1501_),
    .B1_N(_1500_),
    .X(_1503_));
 sky130_fd_sc_hd__xor2_2 _5062_ (.A(_1499_),
    .B(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__a21oi_2 _5063_ (.A1(net106),
    .A2(net177),
    .B1(_1413_),
    .Y(_1505_));
 sky130_fd_sc_hd__a21o_1 _5064_ (.A1(_1411_),
    .A2(_1413_),
    .B1(_1414_),
    .X(_1506_));
 sky130_fd_sc_hd__a21oi_2 _5065_ (.A1(net177),
    .A2(_1506_),
    .B1(_1505_),
    .Y(_1507_));
 sky130_fd_sc_hd__xnor2_2 _5066_ (.A(_1504_),
    .B(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__and2b_1 _5067_ (.A_N(_1508_),
    .B(_1498_),
    .X(_1509_));
 sky130_fd_sc_hd__xnor2_2 _5068_ (.A(_1498_),
    .B(_1508_),
    .Y(_1510_));
 sky130_fd_sc_hd__xnor2_2 _5069_ (.A(_1497_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__nor2_1 _5070_ (.A(_1488_),
    .B(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__xor2_2 _5071_ (.A(_1488_),
    .B(_1511_),
    .X(_1513_));
 sky130_fd_sc_hd__xnor2_2 _5072_ (.A(_1487_),
    .B(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__and2b_1 _5073_ (.A_N(_1514_),
    .B(_1466_),
    .X(_1515_));
 sky130_fd_sc_hd__xnor2_2 _5074_ (.A(_1466_),
    .B(_1514_),
    .Y(_1516_));
 sky130_fd_sc_hd__xnor2_2 _5075_ (.A(_1465_),
    .B(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__nor2_1 _5076_ (.A(_1450_),
    .B(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__xor2_2 _5077_ (.A(_1450_),
    .B(_1517_),
    .X(_1519_));
 sky130_fd_sc_hd__xnor2_1 _5078_ (.A(_1371_),
    .B(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__o21ba_1 _5079_ (.A1(_1433_),
    .A2(_1435_),
    .B1_N(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__or3b_2 _5080_ (.A(_1433_),
    .B(_1435_),
    .C_N(_1520_),
    .X(_1522_));
 sky130_fd_sc_hd__nand2b_1 _5081_ (.A_N(_1521_),
    .B(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__a31o_1 _5082_ (.A1(_1264_),
    .A2(_1347_),
    .A3(_1439_),
    .B1(_1437_),
    .X(_1524_));
 sky130_fd_sc_hd__xnor2_2 _5083_ (.A(_1523_),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nand3_1 _5084_ (.A(_1446_),
    .B(_1449_),
    .C(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__a21o_1 _5085_ (.A1(_1446_),
    .A2(_1449_),
    .B1(_1525_),
    .X(_1527_));
 sky130_fd_sc_hd__a21oi_2 _5086_ (.A1(_1526_),
    .A2(_1527_),
    .B1(net195),
    .Y(_0008_));
 sky130_fd_sc_hd__nor2_1 _5087_ (.A(_1441_),
    .B(_1523_),
    .Y(_1528_));
 sky130_fd_sc_hd__a31o_1 _5088_ (.A1(_1443_),
    .A2(_1444_),
    .A3(_1525_),
    .B1(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__o311a_1 _5089_ (.A1(_1355_),
    .A2(_1357_),
    .A3(_1358_),
    .B1(_1447_),
    .C1(_1525_),
    .X(_1530_));
 sky130_fd_sc_hd__or2_1 _5090_ (.A(_1529_),
    .B(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__a21oi_2 _5091_ (.A1(_1371_),
    .A2(_1519_),
    .B1(_1518_),
    .Y(_1532_));
 sky130_fd_sc_hd__a21o_1 _5092_ (.A1(_1451_),
    .A2(_1462_),
    .B1(_1464_),
    .X(_1533_));
 sky130_fd_sc_hd__a21o_1 _5093_ (.A1(_1465_),
    .A2(_1516_),
    .B1(_1515_),
    .X(_1534_));
 sky130_fd_sc_hd__nand2_2 _5094_ (.A(net135),
    .B(net146),
    .Y(_1535_));
 sky130_fd_sc_hd__and3_2 _5095_ (.A(net135),
    .B(net138),
    .C(net146),
    .X(_1536_));
 sky130_fd_sc_hd__o21ai_1 _5096_ (.A1(net135),
    .A2(net138),
    .B1(net146),
    .Y(_1537_));
 sky130_fd_sc_hd__nand2_1 _5097_ (.A(_1452_),
    .B(_1535_),
    .Y(_1538_));
 sky130_fd_sc_hd__o21a_1 _5098_ (.A1(_1536_),
    .A2(_1537_),
    .B1(_1359_),
    .X(_1539_));
 sky130_fd_sc_hd__nor3_2 _5099_ (.A(_1359_),
    .B(_1536_),
    .C(_1537_),
    .Y(_1540_));
 sky130_fd_sc_hd__nor2_2 _5100_ (.A(_1539_),
    .B(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__or2_2 _5101_ (.A(_1539_),
    .B(_1540_),
    .X(_1542_));
 sky130_fd_sc_hd__o2bb2a_2 _5102_ (.A1_N(net153),
    .A2_N(_1470_),
    .B1(_1471_),
    .B2(_1468_),
    .X(_1543_));
 sky130_fd_sc_hd__nor2_1 _5103_ (.A(_1542_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__xnor2_2 _5104_ (.A(_1541_),
    .B(_1543_),
    .Y(_1545_));
 sky130_fd_sc_hd__a21oi_2 _5105_ (.A1(net144),
    .A2(net146),
    .B1(_1454_),
    .Y(_1546_));
 sky130_fd_sc_hd__nor2_4 _5106_ (.A(_1453_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__xnor2_2 _5107_ (.A(_1545_),
    .B(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__a21o_1 _5108_ (.A1(_1361_),
    .A2(_1457_),
    .B1(_1459_),
    .X(_1549_));
 sky130_fd_sc_hd__or2_1 _5109_ (.A(_1548_),
    .B(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__xnor2_2 _5110_ (.A(_1548_),
    .B(_1549_),
    .Y(_1551_));
 sky130_fd_sc_hd__xor2_2 _5111_ (.A(_1276_),
    .B(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__a21oi_2 _5112_ (.A1(_1467_),
    .A2(_1485_),
    .B1(_1484_),
    .Y(_1553_));
 sky130_fd_sc_hd__nand2b_1 _5113_ (.A_N(_1553_),
    .B(_1552_),
    .Y(_1554_));
 sky130_fd_sc_hd__xnor2_2 _5114_ (.A(_1552_),
    .B(_1553_),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_1364_),
    .B(_1460_),
    .Y(_1556_));
 sky130_fd_sc_hd__inv_2 _5116_ (.A(_1556_),
    .Y(_1557_));
 sky130_fd_sc_hd__or2_1 _5117_ (.A(_1555_),
    .B(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__nand2_1 _5118_ (.A(_1555_),
    .B(_1557_),
    .Y(_1559_));
 sky130_fd_sc_hd__xnor2_1 _5119_ (.A(_1555_),
    .B(_1557_),
    .Y(_1560_));
 sky130_fd_sc_hd__a21oi_2 _5120_ (.A1(_1487_),
    .A2(_1513_),
    .B1(_1512_),
    .Y(_1561_));
 sky130_fd_sc_hd__nand2_1 _5121_ (.A(_1479_),
    .B(_1481_),
    .Y(_1562_));
 sky130_fd_sc_hd__nand2_1 _5122_ (.A(net134),
    .B(net149),
    .Y(_1563_));
 sky130_fd_sc_hd__a22oi_1 _5123_ (.A1(net128),
    .A2(net153),
    .B1(net151),
    .B2(net131),
    .Y(_1564_));
 sky130_fd_sc_hd__and4_1 _5124_ (.A(net128),
    .B(net131),
    .C(net153),
    .D(net151),
    .X(_1565_));
 sky130_fd_sc_hd__nor2_1 _5125_ (.A(_1564_),
    .B(_1565_),
    .Y(_1566_));
 sky130_fd_sc_hd__xnor2_1 _5126_ (.A(_1563_),
    .B(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__a21boi_2 _5127_ (.A1(_1474_),
    .A2(_1475_),
    .B1_N(_1476_),
    .Y(_1568_));
 sky130_fd_sc_hd__a22o_1 _5128_ (.A1(net122),
    .A2(net163),
    .B1(net160),
    .B2(net124),
    .X(_1569_));
 sky130_fd_sc_hd__nand4_1 _5129_ (.A(net122),
    .B(net124),
    .C(net163),
    .D(net160),
    .Y(_1570_));
 sky130_fd_sc_hd__nand4_1 _5130_ (.A(net126),
    .B(net157),
    .C(_1569_),
    .D(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__a22o_1 _5131_ (.A1(net126),
    .A2(net157),
    .B1(_1569_),
    .B2(_1570_),
    .X(_1572_));
 sky130_fd_sc_hd__nand3b_1 _5132_ (.A_N(_1568_),
    .B(_1571_),
    .C(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__a21bo_1 _5133_ (.A1(_1571_),
    .A2(_1572_),
    .B1_N(_1568_),
    .X(_1574_));
 sky130_fd_sc_hd__nand3_1 _5134_ (.A(_1567_),
    .B(_1573_),
    .C(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__a21o_1 _5135_ (.A1(_1573_),
    .A2(_1574_),
    .B1(_1567_),
    .X(_1576_));
 sky130_fd_sc_hd__a21o_1 _5136_ (.A1(_1489_),
    .A2(_1495_),
    .B1(_1494_),
    .X(_1577_));
 sky130_fd_sc_hd__nand3_1 _5137_ (.A(_1575_),
    .B(_1576_),
    .C(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__a21o_1 _5138_ (.A1(_1575_),
    .A2(_1576_),
    .B1(_1577_),
    .X(_1579_));
 sky130_fd_sc_hd__and3_1 _5139_ (.A(_1562_),
    .B(_1578_),
    .C(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__a21oi_1 _5140_ (.A1(_1578_),
    .A2(_1579_),
    .B1(_1562_),
    .Y(_1581_));
 sky130_fd_sc_hd__nor2_1 _5141_ (.A(_1580_),
    .B(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__a21oi_2 _5142_ (.A1(_1497_),
    .A2(_1510_),
    .B1(_1509_),
    .Y(_1583_));
 sky130_fd_sc_hd__nand2_1 _5143_ (.A(_1491_),
    .B(_1492_),
    .Y(_1584_));
 sky130_fd_sc_hd__a22o_1 _5144_ (.A1(net113),
    .A2(net170),
    .B1(net167),
    .B2(net116),
    .X(_1585_));
 sky130_fd_sc_hd__nand4_2 _5145_ (.A(net113),
    .B(net116),
    .C(net170),
    .D(net167),
    .Y(_1586_));
 sky130_fd_sc_hd__nand4_2 _5146_ (.A(net119),
    .B(net165),
    .C(_1585_),
    .D(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__a22o_1 _5147_ (.A1(net119),
    .A2(net165),
    .B1(_1585_),
    .B2(_1586_),
    .X(_1588_));
 sky130_fd_sc_hd__a31o_1 _5148_ (.A1(net113),
    .A2(net171),
    .A3(_1500_),
    .B1(_1502_),
    .X(_1589_));
 sky130_fd_sc_hd__nand3_1 _5149_ (.A(_1587_),
    .B(_1588_),
    .C(_1589_),
    .Y(_1590_));
 sky130_fd_sc_hd__a21o_1 _5150_ (.A1(_1587_),
    .A2(_1588_),
    .B1(_1589_),
    .X(_1591_));
 sky130_fd_sc_hd__nand2_1 _5151_ (.A(_1590_),
    .B(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__xor2_2 _5152_ (.A(_1584_),
    .B(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__and2_1 _5153_ (.A(net177),
    .B(_1414_),
    .X(_1594_));
 sky130_fd_sc_hd__nand2_1 _5154_ (.A(net177),
    .B(_1414_),
    .Y(_1595_));
 sky130_fd_sc_hd__a21o_1 _5155_ (.A1(_1504_),
    .A2(_1507_),
    .B1(_1594_),
    .X(_1596_));
 sky130_fd_sc_hd__a22o_1 _5156_ (.A1(net106),
    .A2(net175),
    .B1(net174),
    .B2(net108),
    .X(_1597_));
 sky130_fd_sc_hd__and3_1 _5157_ (.A(net106),
    .B(net175),
    .C(net174),
    .X(_1598_));
 sky130_fd_sc_hd__nand4_2 _5158_ (.A(net106),
    .B(net108),
    .C(net175),
    .D(net174),
    .Y(_1599_));
 sky130_fd_sc_hd__nand4_1 _5159_ (.A(net110),
    .B(net171),
    .C(_1597_),
    .D(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__a22o_1 _5160_ (.A1(net110),
    .A2(net171),
    .B1(_1597_),
    .B2(_1599_),
    .X(_1601_));
 sky130_fd_sc_hd__nand2_2 _5161_ (.A(_1600_),
    .B(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__or2_4 _5162_ (.A(_1505_),
    .B(_1594_),
    .X(_1603_));
 sky130_fd_sc_hd__xnor2_2 _5163_ (.A(_1602_),
    .B(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__and2b_1 _5164_ (.A_N(_1604_),
    .B(_1596_),
    .X(_1605_));
 sky130_fd_sc_hd__xor2_2 _5165_ (.A(_1596_),
    .B(_1604_),
    .X(_1606_));
 sky130_fd_sc_hd__xnor2_2 _5166_ (.A(_1593_),
    .B(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__nor2_1 _5167_ (.A(_1583_),
    .B(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__xor2_2 _5168_ (.A(_1583_),
    .B(_1607_),
    .X(_1609_));
 sky130_fd_sc_hd__xnor2_1 _5169_ (.A(_1582_),
    .B(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__nor2_1 _5170_ (.A(_1561_),
    .B(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__xor2_1 _5171_ (.A(_1561_),
    .B(_1610_),
    .X(_1612_));
 sky130_fd_sc_hd__xnor2_1 _5172_ (.A(_1560_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(_1534_),
    .B(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__xnor2_1 _5174_ (.A(_1534_),
    .B(_1613_),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2b_1 _5175_ (.A_N(_1615_),
    .B(_1533_),
    .Y(_1616_));
 sky130_fd_sc_hd__xnor2_2 _5176_ (.A(_1533_),
    .B(_1615_),
    .Y(_1617_));
 sky130_fd_sc_hd__and2b_1 _5177_ (.A_N(_1532_),
    .B(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__inv_2 _5178_ (.A(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__xnor2_2 _5179_ (.A(_1532_),
    .B(_1617_),
    .Y(_1620_));
 sky130_fd_sc_hd__a21o_1 _5180_ (.A1(_1437_),
    .A2(_1522_),
    .B1(_1521_),
    .X(_1621_));
 sky130_fd_sc_hd__xnor2_1 _5181_ (.A(_1620_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__inv_2 _5182_ (.A(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__or2_1 _5183_ (.A(_1531_),
    .B(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_1 _5184_ (.A(_1531_),
    .B(_1623_),
    .Y(_1625_));
 sky130_fd_sc_hd__and3_1 _5185_ (.A(net209),
    .B(_1624_),
    .C(_1625_),
    .X(_0009_));
 sky130_fd_sc_hd__and4b_1 _5186_ (.A_N(_1521_),
    .B(_1522_),
    .C(_1620_),
    .D(_1437_),
    .X(_1626_));
 sky130_fd_sc_hd__a21o_1 _5187_ (.A1(_1531_),
    .A2(_1623_),
    .B1(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__nand2_1 _5188_ (.A(_1554_),
    .B(_1559_),
    .Y(_1628_));
 sky130_fd_sc_hd__a31o_1 _5189_ (.A1(_1558_),
    .A2(_1559_),
    .A3(_1612_),
    .B1(_1611_),
    .X(_1629_));
 sky130_fd_sc_hd__o21ai_2 _5190_ (.A1(_1276_),
    .A2(_1551_),
    .B1(_1550_),
    .Y(_1630_));
 sky130_fd_sc_hd__a21oi_2 _5191_ (.A1(_1545_),
    .A2(_1547_),
    .B1(_1544_),
    .Y(_1631_));
 sky130_fd_sc_hd__nor2_2 _5192_ (.A(_1536_),
    .B(_1540_),
    .Y(_1632_));
 sky130_fd_sc_hd__or2_2 _5193_ (.A(_1536_),
    .B(_1540_),
    .X(_1633_));
 sky130_fd_sc_hd__nand2_2 _5194_ (.A(net132),
    .B(net146),
    .Y(_1634_));
 sky130_fd_sc_hd__o21ai_2 _5195_ (.A1(net132),
    .A2(net135),
    .B1(net146),
    .Y(_1635_));
 sky130_fd_sc_hd__and3_1 _5196_ (.A(net132),
    .B(net135),
    .C(net146),
    .X(_1636_));
 sky130_fd_sc_hd__nor2_2 _5197_ (.A(_1635_),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__xnor2_4 _5198_ (.A(_1452_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__a31o_1 _5199_ (.A1(net134),
    .A2(net149),
    .A3(_1566_),
    .B1(_1565_),
    .X(_1639_));
 sky130_fd_sc_hd__and2_1 _5200_ (.A(_1638_),
    .B(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__xor2_1 _5201_ (.A(_1638_),
    .B(_1639_),
    .X(_1641_));
 sky130_fd_sc_hd__and2_1 _5202_ (.A(_1633_),
    .B(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__nor2_1 _5203_ (.A(_1633_),
    .B(_1641_),
    .Y(_1643_));
 sky130_fd_sc_hd__xnor2_1 _5204_ (.A(_1632_),
    .B(_1641_),
    .Y(_1644_));
 sky130_fd_sc_hd__xnor2_2 _5205_ (.A(_1631_),
    .B(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_1363_),
    .B(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__xnor2_2 _5207_ (.A(_1363_),
    .B(_1645_),
    .Y(_1647_));
 sky130_fd_sc_hd__a31o_1 _5208_ (.A1(_1575_),
    .A2(_1576_),
    .A3(_1577_),
    .B1(_1580_),
    .X(_1648_));
 sky130_fd_sc_hd__and2b_1 _5209_ (.A_N(_1647_),
    .B(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__xor2_2 _5210_ (.A(_1647_),
    .B(_1648_),
    .X(_1650_));
 sky130_fd_sc_hd__and2b_1 _5211_ (.A_N(_1650_),
    .B(_1630_),
    .X(_1651_));
 sky130_fd_sc_hd__xnor2_2 _5212_ (.A(_1630_),
    .B(_1650_),
    .Y(_1652_));
 sky130_fd_sc_hd__a21oi_2 _5213_ (.A1(_1582_),
    .A2(_1609_),
    .B1(_1608_),
    .Y(_1653_));
 sky130_fd_sc_hd__and2_1 _5214_ (.A(_1573_),
    .B(_1575_),
    .X(_1654_));
 sky130_fd_sc_hd__a22o_1 _5215_ (.A1(net126),
    .A2(net153),
    .B1(net151),
    .B2(net128),
    .X(_1655_));
 sky130_fd_sc_hd__and4_1 _5216_ (.A(net126),
    .B(net128),
    .C(net153),
    .D(net151),
    .X(_1656_));
 sky130_fd_sc_hd__inv_2 _5217_ (.A(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__and4b_1 _5218_ (.A_N(_1656_),
    .B(net149),
    .C(net131),
    .D(_1655_),
    .X(_1658_));
 sky130_fd_sc_hd__a22oi_1 _5219_ (.A1(net131),
    .A2(net149),
    .B1(_1655_),
    .B2(_1657_),
    .Y(_1659_));
 sky130_fd_sc_hd__nor2_1 _5220_ (.A(_1658_),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__and2_1 _5221_ (.A(_1570_),
    .B(_1571_),
    .X(_1661_));
 sky130_fd_sc_hd__a22oi_1 _5222_ (.A1(net119),
    .A2(net163),
    .B1(net160),
    .B2(net122),
    .Y(_1662_));
 sky130_fd_sc_hd__and4_1 _5223_ (.A(net119),
    .B(net122),
    .C(net163),
    .D(net160),
    .X(_1663_));
 sky130_fd_sc_hd__and4bb_1 _5224_ (.A_N(_1662_),
    .B_N(_1663_),
    .C(net124),
    .D(net157),
    .X(_1664_));
 sky130_fd_sc_hd__o2bb2a_1 _5225_ (.A1_N(net124),
    .A2_N(net157),
    .B1(_1662_),
    .B2(_1663_),
    .X(_1665_));
 sky130_fd_sc_hd__nor2_1 _5226_ (.A(_1664_),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__and2b_1 _5227_ (.A_N(_1661_),
    .B(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__xnor2_2 _5228_ (.A(_1661_),
    .B(_1666_),
    .Y(_1668_));
 sky130_fd_sc_hd__and2_1 _5229_ (.A(_1660_),
    .B(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__xnor2_2 _5230_ (.A(_1660_),
    .B(_1668_),
    .Y(_1670_));
 sky130_fd_sc_hd__a21bo_1 _5231_ (.A1(_1584_),
    .A2(_1591_),
    .B1_N(_1590_),
    .X(_1671_));
 sky130_fd_sc_hd__and2b_1 _5232_ (.A_N(_1670_),
    .B(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__xor2_2 _5233_ (.A(_1670_),
    .B(_1671_),
    .X(_1673_));
 sky130_fd_sc_hd__xor2_2 _5234_ (.A(_1654_),
    .B(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__o21bai_2 _5235_ (.A1(_1593_),
    .A2(_1606_),
    .B1_N(_1605_),
    .Y(_1675_));
 sky130_fd_sc_hd__nand2_2 _5236_ (.A(_1586_),
    .B(_1587_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _5237_ (.A(net116),
    .B(net165),
    .Y(_1677_));
 sky130_fd_sc_hd__a22o_1 _5238_ (.A1(net110),
    .A2(net170),
    .B1(net167),
    .B2(net113),
    .X(_1678_));
 sky130_fd_sc_hd__and3_1 _5239_ (.A(net110),
    .B(net113),
    .C(net167),
    .X(_1679_));
 sky130_fd_sc_hd__a21bo_1 _5240_ (.A1(net170),
    .A2(_1679_),
    .B1_N(_1678_),
    .X(_1680_));
 sky130_fd_sc_hd__xor2_2 _5241_ (.A(_1677_),
    .B(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_1599_),
    .B(_1600_),
    .Y(_1682_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_1681_),
    .B(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__xor2_2 _5244_ (.A(_1681_),
    .B(_1682_),
    .X(_1684_));
 sky130_fd_sc_hd__nand2_1 _5245_ (.A(_1676_),
    .B(_1684_),
    .Y(_1685_));
 sky130_fd_sc_hd__xnor2_2 _5246_ (.A(_1676_),
    .B(_1684_),
    .Y(_1686_));
 sky130_fd_sc_hd__o21ai_2 _5247_ (.A1(_1602_),
    .A2(_1603_),
    .B1(_1595_),
    .Y(_1687_));
 sky130_fd_sc_hd__nand2_1 _5248_ (.A(net108),
    .B(net171),
    .Y(_1688_));
 sky130_fd_sc_hd__o21ai_2 _5249_ (.A1(\ann.weight[3] ),
    .A2(net174),
    .B1(net106),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_2 _5250_ (.A(_1598_),
    .B(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__xnor2_2 _5251_ (.A(_1688_),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__and2b_1 _5252_ (.A_N(_1603_),
    .B(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__xnor2_2 _5253_ (.A(_1603_),
    .B(_1691_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_1 _5254_ (.A(_1687_),
    .B(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__xnor2_2 _5255_ (.A(_1687_),
    .B(_1693_),
    .Y(_1695_));
 sky130_fd_sc_hd__xnor2_2 _5256_ (.A(_1686_),
    .B(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__nand2b_1 _5257_ (.A_N(_1696_),
    .B(_1675_),
    .Y(_1697_));
 sky130_fd_sc_hd__xnor2_2 _5258_ (.A(_1675_),
    .B(_1696_),
    .Y(_1698_));
 sky130_fd_sc_hd__xnor2_2 _5259_ (.A(_1674_),
    .B(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_1 _5260_ (.A(_1653_),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__xor2_2 _5261_ (.A(_1653_),
    .B(_1699_),
    .X(_1701_));
 sky130_fd_sc_hd__xor2_1 _5262_ (.A(_1652_),
    .B(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__nand2_1 _5263_ (.A(_1629_),
    .B(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__xor2_1 _5264_ (.A(_1629_),
    .B(_1702_),
    .X(_1704_));
 sky130_fd_sc_hd__xnor2_1 _5265_ (.A(_1628_),
    .B(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__a21oi_2 _5266_ (.A1(_1614_),
    .A2(_1616_),
    .B1(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__inv_2 _5267_ (.A(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__and3_1 _5268_ (.A(_1614_),
    .B(_1616_),
    .C(_1705_),
    .X(_1708_));
 sky130_fd_sc_hd__or2_1 _5269_ (.A(_1706_),
    .B(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__nand2_1 _5270_ (.A(_1521_),
    .B(_1620_),
    .Y(_1710_));
 sky130_fd_sc_hd__a21o_1 _5271_ (.A1(_1521_),
    .A2(_1620_),
    .B1(_1618_),
    .X(_1711_));
 sky130_fd_sc_hd__xnor2_1 _5272_ (.A(_1709_),
    .B(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__xnor2_1 _5273_ (.A(_1627_),
    .B(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__nor2_1 _5274_ (.A(net194),
    .B(_1713_),
    .Y(_0010_));
 sky130_fd_sc_hd__and2b_1 _5275_ (.A_N(_1622_),
    .B(_1712_),
    .X(_1714_));
 sky130_fd_sc_hd__nor2_1 _5276_ (.A(_1709_),
    .B(_1710_),
    .Y(_1715_));
 sky130_fd_sc_hd__a221o_1 _5277_ (.A1(_1626_),
    .A2(_1712_),
    .B1(_1714_),
    .B2(_1529_),
    .C1(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__a21oi_2 _5278_ (.A1(_1530_),
    .A2(_1714_),
    .B1(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hd__a21bo_1 _5279_ (.A1(_1628_),
    .A2(_1704_),
    .B1_N(_1703_),
    .X(_1718_));
 sky130_fd_sc_hd__nor2_1 _5280_ (.A(_1649_),
    .B(_1651_),
    .Y(_1719_));
 sky130_fd_sc_hd__a21oi_2 _5281_ (.A1(_1652_),
    .A2(_1701_),
    .B1(_1700_),
    .Y(_1720_));
 sky130_fd_sc_hd__o31a_1 _5282_ (.A1(_1631_),
    .A2(_1642_),
    .A3(_1643_),
    .B1(_1646_),
    .X(_1721_));
 sky130_fd_sc_hd__and4_2 _5283_ (.A(net138),
    .B(net142),
    .C(net144),
    .D(net146),
    .X(_1722_));
 sky130_fd_sc_hd__o21bai_4 _5284_ (.A1(_1360_),
    .A2(_1456_),
    .B1_N(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__o21ba_4 _5285_ (.A1(_1452_),
    .A2(_1635_),
    .B1_N(_1636_),
    .X(_1724_));
 sky130_fd_sc_hd__inv_2 _5286_ (.A(_1724_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_2 _5287_ (.A(net129),
    .B(net147),
    .Y(_1726_));
 sky130_fd_sc_hd__o21ai_2 _5288_ (.A1(net129),
    .A2(net132),
    .B1(net146),
    .Y(_1727_));
 sky130_fd_sc_hd__and3_1 _5289_ (.A(net129),
    .B(net132),
    .C(net146),
    .X(_1728_));
 sky130_fd_sc_hd__nor2_2 _5290_ (.A(_1727_),
    .B(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hd__xnor2_4 _5291_ (.A(_1535_),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__nor2_1 _5292_ (.A(_1656_),
    .B(_1658_),
    .Y(_1731_));
 sky130_fd_sc_hd__and2b_1 _5293_ (.A_N(_1731_),
    .B(_1730_),
    .X(_1732_));
 sky130_fd_sc_hd__xnor2_1 _5294_ (.A(_1730_),
    .B(_1731_),
    .Y(_1733_));
 sky130_fd_sc_hd__and2_1 _5295_ (.A(_1725_),
    .B(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__xnor2_1 _5296_ (.A(_1724_),
    .B(_1733_),
    .Y(_1735_));
 sky130_fd_sc_hd__o21ai_2 _5297_ (.A1(_1640_),
    .A2(_1642_),
    .B1(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__or3_1 _5298_ (.A(_1640_),
    .B(_1642_),
    .C(_1735_),
    .X(_1737_));
 sky130_fd_sc_hd__nand2_1 _5299_ (.A(_1736_),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__or2_1 _5300_ (.A(_1723_),
    .B(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__xor2_2 _5301_ (.A(_1723_),
    .B(_1738_),
    .X(_1740_));
 sky130_fd_sc_hd__o21ba_1 _5302_ (.A1(_1654_),
    .A2(_1673_),
    .B1_N(_1672_),
    .X(_1741_));
 sky130_fd_sc_hd__and2b_1 _5303_ (.A_N(_1741_),
    .B(_1740_),
    .X(_1742_));
 sky130_fd_sc_hd__xnor2_2 _5304_ (.A(_1740_),
    .B(_1741_),
    .Y(_1743_));
 sky130_fd_sc_hd__and2b_1 _5305_ (.A_N(_1721_),
    .B(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__xnor2_2 _5306_ (.A(_1721_),
    .B(_1743_),
    .Y(_1745_));
 sky130_fd_sc_hd__a21bo_1 _5307_ (.A1(_1674_),
    .A2(_1698_),
    .B1_N(_1697_),
    .X(_1746_));
 sky130_fd_sc_hd__a22o_1 _5308_ (.A1(net124),
    .A2(net153),
    .B1(net151),
    .B2(net126),
    .X(_1747_));
 sky130_fd_sc_hd__and4_1 _5309_ (.A(net124),
    .B(net126),
    .C(net153),
    .D(net151),
    .X(_1748_));
 sky130_fd_sc_hd__inv_2 _5310_ (.A(_1748_),
    .Y(_1749_));
 sky130_fd_sc_hd__a22oi_1 _5311_ (.A1(net128),
    .A2(net149),
    .B1(_1747_),
    .B2(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__and4b_1 _5312_ (.A_N(_1748_),
    .B(net149),
    .C(net128),
    .D(_1747_),
    .X(_1751_));
 sky130_fd_sc_hd__nor2_1 _5313_ (.A(_1750_),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__or2_1 _5314_ (.A(_1663_),
    .B(_1664_),
    .X(_1753_));
 sky130_fd_sc_hd__a22oi_1 _5315_ (.A1(net116),
    .A2(net163),
    .B1(net160),
    .B2(net119),
    .Y(_1754_));
 sky130_fd_sc_hd__and4_1 _5316_ (.A(net116),
    .B(net119),
    .C(net163),
    .D(net160),
    .X(_1755_));
 sky130_fd_sc_hd__o2bb2a_1 _5317_ (.A1_N(net122),
    .A2_N(net157),
    .B1(_1754_),
    .B2(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__and4bb_1 _5318_ (.A_N(_1754_),
    .B_N(_1755_),
    .C(net122),
    .D(net157),
    .X(_1757_));
 sky130_fd_sc_hd__nor2_1 _5319_ (.A(_1756_),
    .B(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__and2_1 _5320_ (.A(_1753_),
    .B(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__xor2_1 _5321_ (.A(_1753_),
    .B(_1758_),
    .X(_1760_));
 sky130_fd_sc_hd__and2_1 _5322_ (.A(_1752_),
    .B(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__xnor2_1 _5323_ (.A(_1752_),
    .B(_1760_),
    .Y(_1762_));
 sky130_fd_sc_hd__a21o_1 _5324_ (.A1(_1683_),
    .A2(_1685_),
    .B1(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__nand3_1 _5325_ (.A(_1683_),
    .B(_1685_),
    .C(_1762_),
    .Y(_1764_));
 sky130_fd_sc_hd__o211ai_2 _5326_ (.A1(_1667_),
    .A2(_1669_),
    .B1(_1763_),
    .C1(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__a211o_1 _5327_ (.A1(_1763_),
    .A2(_1764_),
    .B1(_1667_),
    .C1(_1669_),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_1 _5328_ (.A(_1765_),
    .B(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__o21ai_2 _5329_ (.A1(_1686_),
    .A2(_1695_),
    .B1(_1694_),
    .Y(_1768_));
 sky130_fd_sc_hd__a32o_1 _5330_ (.A1(net116),
    .A2(net165),
    .A3(_1678_),
    .B1(_1679_),
    .B2(net170),
    .X(_1769_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(net108),
    .A2(net170),
    .B1(net167),
    .B2(net110),
    .X(_1770_));
 sky130_fd_sc_hd__inv_2 _5332_ (.A(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__and4_1 _5333_ (.A(net108),
    .B(net110),
    .C(net170),
    .D(net167),
    .X(_1772_));
 sky130_fd_sc_hd__o2bb2a_1 _5334_ (.A1_N(net113),
    .A2_N(net165),
    .B1(_1771_),
    .B2(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__and4b_1 _5335_ (.A_N(_1772_),
    .B(net165),
    .C(net113),
    .D(_1770_),
    .X(_1774_));
 sky130_fd_sc_hd__nor2_1 _5336_ (.A(_1773_),
    .B(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__o21ba_1 _5337_ (.A1(_1688_),
    .A2(_1689_),
    .B1_N(_1598_),
    .X(_1776_));
 sky130_fd_sc_hd__or3_1 _5338_ (.A(_1773_),
    .B(_1774_),
    .C(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__xnor2_2 _5339_ (.A(_1775_),
    .B(_1776_),
    .Y(_1778_));
 sky130_fd_sc_hd__nand2_1 _5340_ (.A(_1769_),
    .B(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__xor2_2 _5341_ (.A(_1769_),
    .B(_1778_),
    .X(_1780_));
 sky130_fd_sc_hd__nand2_1 _5342_ (.A(net106),
    .B(net171),
    .Y(_1781_));
 sky130_fd_sc_hd__xor2_2 _5343_ (.A(_1690_),
    .B(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__xor2_1 _5344_ (.A(_1603_),
    .B(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__o21ai_1 _5345_ (.A1(_1594_),
    .A2(_1692_),
    .B1(_1783_),
    .Y(_1784_));
 sky130_fd_sc_hd__or3_1 _5346_ (.A(_1594_),
    .B(_1692_),
    .C(_1783_),
    .X(_1785_));
 sky130_fd_sc_hd__and2_1 _5347_ (.A(_1784_),
    .B(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__nand2_1 _5348_ (.A(_1780_),
    .B(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__xnor2_2 _5349_ (.A(_1780_),
    .B(_1786_),
    .Y(_1788_));
 sky130_fd_sc_hd__nand2b_1 _5350_ (.A_N(_1788_),
    .B(_1768_),
    .Y(_1789_));
 sky130_fd_sc_hd__xnor2_2 _5351_ (.A(_1768_),
    .B(_1788_),
    .Y(_1790_));
 sky130_fd_sc_hd__nand2b_1 _5352_ (.A_N(_1767_),
    .B(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__xnor2_2 _5353_ (.A(_1767_),
    .B(_1790_),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _5354_ (.A(_1746_),
    .B(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__or2_1 _5355_ (.A(_1746_),
    .B(_1792_),
    .X(_1794_));
 sky130_fd_sc_hd__xnor2_1 _5356_ (.A(_1746_),
    .B(_1792_),
    .Y(_1795_));
 sky130_fd_sc_hd__nand3_1 _5357_ (.A(_1745_),
    .B(_1793_),
    .C(_1794_),
    .Y(_1796_));
 sky130_fd_sc_hd__xnor2_2 _5358_ (.A(_1745_),
    .B(_1795_),
    .Y(_1797_));
 sky130_fd_sc_hd__and2b_1 _5359_ (.A_N(_1720_),
    .B(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__xnor2_2 _5360_ (.A(_1720_),
    .B(_1797_),
    .Y(_1799_));
 sky130_fd_sc_hd__and2b_1 _5361_ (.A_N(_1719_),
    .B(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__xnor2_2 _5362_ (.A(_1719_),
    .B(_1799_),
    .Y(_1801_));
 sky130_fd_sc_hd__and2_1 _5363_ (.A(_1718_),
    .B(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__xnor2_2 _5364_ (.A(_1718_),
    .B(_1801_),
    .Y(_1803_));
 sky130_fd_sc_hd__nor2_1 _5365_ (.A(_1619_),
    .B(_1709_),
    .Y(_1804_));
 sky130_fd_sc_hd__nor2_1 _5366_ (.A(_1706_),
    .B(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__xnor2_2 _5367_ (.A(_1803_),
    .B(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__o21ai_1 _5368_ (.A1(_1717_),
    .A2(_1806_),
    .B1(net209),
    .Y(_1807_));
 sky130_fd_sc_hd__a21oi_1 _5369_ (.A1(_1717_),
    .A2(_1806_),
    .B1(_1807_),
    .Y(_0012_));
 sky130_fd_sc_hd__and2b_1 _5370_ (.A_N(_1803_),
    .B(_1804_),
    .X(_1808_));
 sky130_fd_sc_hd__o21bai_1 _5371_ (.A1(_1717_),
    .A2(_1806_),
    .B1_N(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__nor2_1 _5372_ (.A(_1798_),
    .B(_1800_),
    .Y(_1810_));
 sky130_fd_sc_hd__or2_1 _5373_ (.A(_1798_),
    .B(_1800_),
    .X(_1811_));
 sky130_fd_sc_hd__or2_1 _5374_ (.A(_1742_),
    .B(_1744_),
    .X(_1812_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(_1722_),
    .B(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__or2_1 _5376_ (.A(_1722_),
    .B(_1812_),
    .X(_1814_));
 sky130_fd_sc_hd__nand2_1 _5377_ (.A(_1813_),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(_1541_),
    .B(_1547_),
    .Y(_1816_));
 sky130_fd_sc_hd__or2_1 _5379_ (.A(_1541_),
    .B(_1547_),
    .X(_1817_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(_1816_),
    .B(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__or2_1 _5381_ (.A(_1276_),
    .B(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__nand2_1 _5382_ (.A(_1276_),
    .B(_1818_),
    .Y(_1820_));
 sky130_fd_sc_hd__and2_2 _5383_ (.A(_1819_),
    .B(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__o21ba_4 _5384_ (.A1(_1535_),
    .A2(_1727_),
    .B1_N(_1728_),
    .X(_1822_));
 sky130_fd_sc_hd__nand2_2 _5385_ (.A(net127),
    .B(net147),
    .Y(_1823_));
 sky130_fd_sc_hd__o21ai_1 _5386_ (.A1(net127),
    .A2(net129),
    .B1(net146),
    .Y(_1824_));
 sky130_fd_sc_hd__and3_1 _5387_ (.A(net127),
    .B(net129),
    .C(net146),
    .X(_1825_));
 sky130_fd_sc_hd__nor2_2 _5388_ (.A(_1824_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__xnor2_4 _5389_ (.A(_1634_),
    .B(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__nor2_1 _5390_ (.A(_1748_),
    .B(_1751_),
    .Y(_1828_));
 sky130_fd_sc_hd__and2b_1 _5391_ (.A_N(_1828_),
    .B(_1827_),
    .X(_1829_));
 sky130_fd_sc_hd__xnor2_1 _5392_ (.A(_1827_),
    .B(_1828_),
    .Y(_1830_));
 sky130_fd_sc_hd__and2b_1 _5393_ (.A_N(_1822_),
    .B(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__xnor2_1 _5394_ (.A(_1822_),
    .B(_1830_),
    .Y(_1832_));
 sky130_fd_sc_hd__o21ai_2 _5395_ (.A1(_1732_),
    .A2(_1734_),
    .B1(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__or3_1 _5396_ (.A(_1732_),
    .B(_1734_),
    .C(_1832_),
    .X(_1834_));
 sky130_fd_sc_hd__and2_1 _5397_ (.A(_1833_),
    .B(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__nand2_1 _5398_ (.A(_1821_),
    .B(_1835_),
    .Y(_1836_));
 sky130_fd_sc_hd__xnor2_1 _5399_ (.A(_1821_),
    .B(_1835_),
    .Y(_1837_));
 sky130_fd_sc_hd__a21oi_2 _5400_ (.A1(_1763_),
    .A2(_1765_),
    .B1(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__and3_1 _5401_ (.A(_1763_),
    .B(_1765_),
    .C(_1837_),
    .X(_1839_));
 sky130_fd_sc_hd__a211oi_2 _5402_ (.A1(_1736_),
    .A2(_1739_),
    .B1(_1838_),
    .C1(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__o211a_1 _5403_ (.A1(_1838_),
    .A2(_1839_),
    .B1(_1736_),
    .C1(_1739_),
    .X(_1841_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(net126),
    .B(net149),
    .Y(_1842_));
 sky130_fd_sc_hd__a22o_1 _5405_ (.A1(net122),
    .A2(net153),
    .B1(net151),
    .B2(net124),
    .X(_1843_));
 sky130_fd_sc_hd__and3_1 _5406_ (.A(net122),
    .B(net124),
    .C(net151),
    .X(_1844_));
 sky130_fd_sc_hd__a21bo_1 _5407_ (.A1(net153),
    .A2(_1844_),
    .B1_N(_1843_),
    .X(_1845_));
 sky130_fd_sc_hd__xor2_1 _5408_ (.A(_1842_),
    .B(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__or2_1 _5409_ (.A(_1755_),
    .B(_1757_),
    .X(_1847_));
 sky130_fd_sc_hd__a22o_1 _5410_ (.A1(net113),
    .A2(net161),
    .B1(net158),
    .B2(net115),
    .X(_1848_));
 sky130_fd_sc_hd__and4_1 _5411_ (.A(net113),
    .B(net115),
    .C(net161),
    .D(net158),
    .X(_1849_));
 sky130_fd_sc_hd__inv_2 _5412_ (.A(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__a22oi_1 _5413_ (.A1(net118),
    .A2(net157),
    .B1(_1848_),
    .B2(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__and4_1 _5414_ (.A(net118),
    .B(net157),
    .C(_1848_),
    .D(_1850_),
    .X(_1852_));
 sky130_fd_sc_hd__nor2_1 _5415_ (.A(_1851_),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__and2_1 _5416_ (.A(_1847_),
    .B(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__xor2_1 _5417_ (.A(_1847_),
    .B(_1853_),
    .X(_1855_));
 sky130_fd_sc_hd__and2_1 _5418_ (.A(_1846_),
    .B(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__xnor2_1 _5419_ (.A(_1846_),
    .B(_1855_),
    .Y(_1857_));
 sky130_fd_sc_hd__a21o_1 _5420_ (.A1(_1777_),
    .A2(_1779_),
    .B1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__nand3_1 _5421_ (.A(_1777_),
    .B(_1779_),
    .C(_1857_),
    .Y(_1859_));
 sky130_fd_sc_hd__o211a_1 _5422_ (.A1(_1759_),
    .A2(_1761_),
    .B1(_1858_),
    .C1(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__inv_2 _5423_ (.A(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__a211oi_1 _5424_ (.A1(_1858_),
    .A2(_1859_),
    .B1(_1759_),
    .C1(_1761_),
    .Y(_1862_));
 sky130_fd_sc_hd__or2_1 _5425_ (.A(_1860_),
    .B(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__nand2_1 _5426_ (.A(_1784_),
    .B(_1787_),
    .Y(_1864_));
 sky130_fd_sc_hd__or2_1 _5427_ (.A(_1772_),
    .B(_1774_),
    .X(_1865_));
 sky130_fd_sc_hd__a22oi_1 _5428_ (.A1(net106),
    .A2(net170),
    .B1(net167),
    .B2(net108),
    .Y(_1866_));
 sky130_fd_sc_hd__and4_1 _5429_ (.A(net106),
    .B(net108),
    .C(net170),
    .D(net167),
    .X(_1867_));
 sky130_fd_sc_hd__nor2_1 _5430_ (.A(_1866_),
    .B(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__a21oi_1 _5431_ (.A1(net110),
    .A2(net165),
    .B1(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__and3_1 _5432_ (.A(net110),
    .B(net165),
    .C(_1868_),
    .X(_1870_));
 sky130_fd_sc_hd__or2_1 _5433_ (.A(_1869_),
    .B(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__o21ba_4 _5434_ (.A1(_1689_),
    .A2(_1781_),
    .B1_N(_1598_),
    .X(_1872_));
 sky130_fd_sc_hd__or2_1 _5435_ (.A(_1871_),
    .B(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__xor2_1 _5436_ (.A(_1871_),
    .B(_1872_),
    .X(_1874_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_1865_),
    .B(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__xnor2_1 _5438_ (.A(_1865_),
    .B(_1874_),
    .Y(_1876_));
 sky130_fd_sc_hd__nor2_1 _5439_ (.A(_1595_),
    .B(_1782_),
    .Y(_1877_));
 sky130_fd_sc_hd__inv_2 _5440_ (.A(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__and2_2 _5441_ (.A(_1505_),
    .B(_1782_),
    .X(_1879_));
 sky130_fd_sc_hd__nor2_2 _5442_ (.A(_1877_),
    .B(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__xor2_1 _5443_ (.A(_1876_),
    .B(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__a21o_1 _5444_ (.A1(_1784_),
    .A2(_1787_),
    .B1(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__xor2_1 _5445_ (.A(_1864_),
    .B(_1881_),
    .X(_1883_));
 sky130_fd_sc_hd__or2_1 _5446_ (.A(_1863_),
    .B(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__xnor2_1 _5447_ (.A(_1863_),
    .B(_1883_),
    .Y(_1885_));
 sky130_fd_sc_hd__a21o_1 _5448_ (.A1(_1789_),
    .A2(_1791_),
    .B1(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__nand3_1 _5449_ (.A(_1789_),
    .B(_1791_),
    .C(_1885_),
    .Y(_1887_));
 sky130_fd_sc_hd__and4bb_1 _5450_ (.A_N(_1840_),
    .B_N(_1841_),
    .C(_1886_),
    .D(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__or4bb_1 _5451_ (.A(_1840_),
    .B(_1841_),
    .C_N(_1886_),
    .D_N(_1887_),
    .X(_1889_));
 sky130_fd_sc_hd__a2bb2oi_1 _5452_ (.A1_N(_1840_),
    .A2_N(_1841_),
    .B1(_1886_),
    .B2(_1887_),
    .Y(_1890_));
 sky130_fd_sc_hd__a211oi_1 _5453_ (.A1(_1793_),
    .A2(_1796_),
    .B1(_1888_),
    .C1(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__o211a_1 _5454_ (.A1(_1888_),
    .A2(_1890_),
    .B1(_1793_),
    .C1(_1796_),
    .X(_1892_));
 sky130_fd_sc_hd__or3_1 _5455_ (.A(_1815_),
    .B(_1891_),
    .C(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__o21ai_1 _5456_ (.A1(_1891_),
    .A2(_1892_),
    .B1(_1815_),
    .Y(_1894_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(_1893_),
    .B(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__xnor2_2 _5458_ (.A(_1811_),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__nor2_1 _5459_ (.A(_1707_),
    .B(_1803_),
    .Y(_1897_));
 sky130_fd_sc_hd__nor2_1 _5460_ (.A(_1802_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__xnor2_1 _5461_ (.A(_1896_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__xnor2_1 _5462_ (.A(_1809_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__nor2_1 _5463_ (.A(net194),
    .B(_1900_),
    .Y(_0013_));
 sky130_fd_sc_hd__a22oi_1 _5464_ (.A1(_1896_),
    .A2(_1897_),
    .B1(_1899_),
    .B2(_1808_),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2b_1 _5465_ (.A_N(_1806_),
    .B(_1899_),
    .Y(_1902_));
 sky130_fd_sc_hd__o21ai_1 _5466_ (.A1(_1717_),
    .A2(_1902_),
    .B1(_1901_),
    .Y(_1903_));
 sky130_fd_sc_hd__o21bai_1 _5467_ (.A1(_1815_),
    .A2(_1892_),
    .B1_N(_1891_),
    .Y(_1904_));
 sky130_fd_sc_hd__nor2_1 _5468_ (.A(_1838_),
    .B(_1840_),
    .Y(_1905_));
 sky130_fd_sc_hd__a21o_1 _5469_ (.A1(_1816_),
    .A2(_1819_),
    .B1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__nand3_1 _5470_ (.A(_1816_),
    .B(_1819_),
    .C(_1905_),
    .Y(_1907_));
 sky130_fd_sc_hd__nand2_1 _5471_ (.A(_1906_),
    .B(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__and2_1 _5472_ (.A(_1633_),
    .B(_1638_),
    .X(_1909_));
 sky130_fd_sc_hd__nor2_1 _5473_ (.A(_1633_),
    .B(_1638_),
    .Y(_1910_));
 sky130_fd_sc_hd__nor2_4 _5474_ (.A(_1909_),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__xnor2_1 _5475_ (.A(_1363_),
    .B(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__o21ba_2 _5476_ (.A1(_1634_),
    .A2(_1824_),
    .B1_N(_1825_),
    .X(_1913_));
 sky130_fd_sc_hd__nand2_2 _5477_ (.A(net125),
    .B(net148),
    .Y(_1914_));
 sky130_fd_sc_hd__o21ai_1 _5478_ (.A1(net125),
    .A2(net127),
    .B1(net147),
    .Y(_1915_));
 sky130_fd_sc_hd__and3_1 _5479_ (.A(net125),
    .B(net127),
    .C(net147),
    .X(_1916_));
 sky130_fd_sc_hd__nor2_2 _5480_ (.A(_1915_),
    .B(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__xnor2_4 _5481_ (.A(_1726_),
    .B(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__a32o_1 _5482_ (.A1(net126),
    .A2(net149),
    .A3(_1843_),
    .B1(_1844_),
    .B2(net153),
    .X(_1919_));
 sky130_fd_sc_hd__and2_1 _5483_ (.A(_1918_),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__nor2_1 _5484_ (.A(_1918_),
    .B(_1919_),
    .Y(_1921_));
 sky130_fd_sc_hd__nor2_1 _5485_ (.A(_1920_),
    .B(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__xnor2_1 _5486_ (.A(_1913_),
    .B(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__o21ai_1 _5487_ (.A1(_1829_),
    .A2(_1831_),
    .B1(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__or3_1 _5488_ (.A(_1829_),
    .B(_1831_),
    .C(_1923_),
    .X(_1925_));
 sky130_fd_sc_hd__nand2_1 _5489_ (.A(_1924_),
    .B(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__or2_1 _5490_ (.A(_1912_),
    .B(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__xnor2_1 _5491_ (.A(_1912_),
    .B(_1926_),
    .Y(_1928_));
 sky130_fd_sc_hd__a21oi_2 _5492_ (.A1(_1858_),
    .A2(_1861_),
    .B1(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__and3_1 _5493_ (.A(_1858_),
    .B(_1861_),
    .C(_1928_),
    .X(_1930_));
 sky130_fd_sc_hd__a211oi_2 _5494_ (.A1(_1833_),
    .A2(_1836_),
    .B1(_1929_),
    .C1(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__o211a_1 _5495_ (.A1(_1929_),
    .A2(_1930_),
    .B1(_1833_),
    .C1(_1836_),
    .X(_1932_));
 sky130_fd_sc_hd__nand2_1 _5496_ (.A(net123),
    .B(net149),
    .Y(_1933_));
 sky130_fd_sc_hd__a22o_1 _5497_ (.A1(net118),
    .A2(net153),
    .B1(net151),
    .B2(net121),
    .X(_1934_));
 sky130_fd_sc_hd__and3_1 _5498_ (.A(net118),
    .B(net121),
    .C(net151),
    .X(_1935_));
 sky130_fd_sc_hd__a21bo_1 _5499_ (.A1(net153),
    .A2(_1935_),
    .B1_N(_1934_),
    .X(_1936_));
 sky130_fd_sc_hd__xor2_1 _5500_ (.A(_1933_),
    .B(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__nor2_1 _5501_ (.A(_1849_),
    .B(_1852_),
    .Y(_1938_));
 sky130_fd_sc_hd__a22o_1 _5502_ (.A1(\ann.in_ff[2][13] ),
    .A2(net161),
    .B1(net158),
    .B2(net112),
    .X(_1939_));
 sky130_fd_sc_hd__and4_1 _5503_ (.A(\ann.in_ff[2][13] ),
    .B(net112),
    .C(net161),
    .D(net158),
    .X(_1940_));
 sky130_fd_sc_hd__inv_2 _5504_ (.A(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__a22oi_1 _5505_ (.A1(net115),
    .A2(net156),
    .B1(_1939_),
    .B2(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__and4b_1 _5506_ (.A_N(_1940_),
    .B(net156),
    .C(net115),
    .D(_1939_),
    .X(_1943_));
 sky130_fd_sc_hd__nor2_1 _5507_ (.A(_1942_),
    .B(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__and2b_1 _5508_ (.A_N(_1938_),
    .B(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__xnor2_1 _5509_ (.A(_1938_),
    .B(_1944_),
    .Y(_1946_));
 sky130_fd_sc_hd__xnor2_1 _5510_ (.A(_1937_),
    .B(_1946_),
    .Y(_1947_));
 sky130_fd_sc_hd__a21o_1 _5511_ (.A1(_1873_),
    .A2(_1875_),
    .B1(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__nand3_1 _5512_ (.A(_1873_),
    .B(_1875_),
    .C(_1947_),
    .Y(_1949_));
 sky130_fd_sc_hd__o211a_1 _5513_ (.A1(_1854_),
    .A2(_1856_),
    .B1(_1948_),
    .C1(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__inv_2 _5514_ (.A(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hd__a211oi_1 _5515_ (.A1(_1948_),
    .A2(_1949_),
    .B1(_1854_),
    .C1(_1856_),
    .Y(_1952_));
 sky130_fd_sc_hd__o21ai_1 _5516_ (.A1(_1876_),
    .A2(_1879_),
    .B1(_1878_),
    .Y(_1953_));
 sky130_fd_sc_hd__or2_1 _5517_ (.A(_1867_),
    .B(_1870_),
    .X(_1954_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(\ann.in_ff[2][14] ),
    .B(net164),
    .Y(_1955_));
 sky130_fd_sc_hd__and3_1 _5519_ (.A(net105),
    .B(net168),
    .C(net166),
    .X(_1956_));
 sky130_fd_sc_hd__o21ai_2 _5520_ (.A1(net168),
    .A2(net166),
    .B1(net105),
    .Y(_1957_));
 sky130_fd_sc_hd__nor2_4 _5521_ (.A(_1956_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__xnor2_2 _5522_ (.A(_1955_),
    .B(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nand2b_1 _5523_ (.A_N(_1872_),
    .B(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__xnor2_1 _5524_ (.A(_1872_),
    .B(_1959_),
    .Y(_1961_));
 sky130_fd_sc_hd__nand2_1 _5525_ (.A(_1954_),
    .B(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__xnor2_1 _5526_ (.A(_1954_),
    .B(_1961_),
    .Y(_1963_));
 sky130_fd_sc_hd__xnor2_1 _5527_ (.A(_1880_),
    .B(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__and2_1 _5528_ (.A(_1953_),
    .B(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__nor2_1 _5529_ (.A(_1953_),
    .B(_1964_),
    .Y(_1966_));
 sky130_fd_sc_hd__or2_1 _5530_ (.A(_1965_),
    .B(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__nor3_2 _5531_ (.A(_1950_),
    .B(_1952_),
    .C(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__o21a_1 _5532_ (.A1(_1950_),
    .A2(_1952_),
    .B1(_1967_),
    .X(_1969_));
 sky130_fd_sc_hd__a211oi_4 _5533_ (.A1(_1882_),
    .A2(_1884_),
    .B1(_1968_),
    .C1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__o211a_1 _5534_ (.A1(_1968_),
    .A2(_1969_),
    .B1(_1882_),
    .C1(_1884_),
    .X(_1971_));
 sky130_fd_sc_hd__nor4_2 _5535_ (.A(_1931_),
    .B(_1932_),
    .C(_1970_),
    .D(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__o22a_1 _5536_ (.A1(_1931_),
    .A2(_1932_),
    .B1(_1970_),
    .B2(_1971_),
    .X(_1973_));
 sky130_fd_sc_hd__a211oi_2 _5537_ (.A1(_1886_),
    .A2(_1889_),
    .B1(net57),
    .C1(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__o211a_1 _5538_ (.A1(net57),
    .A2(_1973_),
    .B1(_1886_),
    .C1(_1889_),
    .X(_1975_));
 sky130_fd_sc_hd__nor3_1 _5539_ (.A(_1908_),
    .B(_1974_),
    .C(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__o21a_1 _5540_ (.A1(_1974_),
    .A2(_1975_),
    .B1(_1908_),
    .X(_1977_));
 sky130_fd_sc_hd__or2_1 _5541_ (.A(_1976_),
    .B(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__and2b_1 _5542_ (.A_N(_1978_),
    .B(_1904_),
    .X(_1979_));
 sky130_fd_sc_hd__xnor2_1 _5543_ (.A(_1904_),
    .B(_1978_),
    .Y(_1980_));
 sky130_fd_sc_hd__xor2_1 _5544_ (.A(_1813_),
    .B(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__nand2_1 _5545_ (.A(_1802_),
    .B(_1896_),
    .Y(_1982_));
 sky130_fd_sc_hd__o21ai_1 _5546_ (.A1(_1810_),
    .A2(_1895_),
    .B1(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__or3b_1 _5547_ (.A(_1895_),
    .B(_1981_),
    .C_N(_1811_),
    .X(_1984_));
 sky130_fd_sc_hd__xnor2_1 _5548_ (.A(_1981_),
    .B(_1983_),
    .Y(_1985_));
 sky130_fd_sc_hd__a21oi_1 _5549_ (.A1(_1903_),
    .A2(_1985_),
    .B1(net195),
    .Y(_1986_));
 sky130_fd_sc_hd__o21a_1 _5550_ (.A1(_1903_),
    .A2(_1985_),
    .B1(_1986_),
    .X(_0014_));
 sky130_fd_sc_hd__a31o_1 _5551_ (.A1(_1722_),
    .A2(_1812_),
    .A3(_1980_),
    .B1(_1979_),
    .X(_1987_));
 sky130_fd_sc_hd__or2_1 _5552_ (.A(_1929_),
    .B(_1931_),
    .X(_1988_));
 sky130_fd_sc_hd__nand2_1 _5553_ (.A(_1360_),
    .B(_1909_),
    .Y(_1989_));
 sky130_fd_sc_hd__or2_1 _5554_ (.A(_1360_),
    .B(_1909_),
    .X(_1990_));
 sky130_fd_sc_hd__a22o_1 _5555_ (.A1(_1363_),
    .A2(_1911_),
    .B1(_1989_),
    .B2(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__nand2_1 _5556_ (.A(_1988_),
    .B(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__xnor2_1 _5557_ (.A(_1988_),
    .B(_1991_),
    .Y(_1993_));
 sky130_fd_sc_hd__xnor2_1 _5558_ (.A(_1724_),
    .B(_1730_),
    .Y(_1994_));
 sky130_fd_sc_hd__and2_1 _5559_ (.A(_1456_),
    .B(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__nor2_1 _5560_ (.A(_1456_),
    .B(_1994_),
    .Y(_1996_));
 sky130_fd_sc_hd__or2_1 _5561_ (.A(_1995_),
    .B(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__o21bai_1 _5562_ (.A1(_1913_),
    .A2(_1921_),
    .B1_N(_1920_),
    .Y(_1998_));
 sky130_fd_sc_hd__o21ba_2 _5563_ (.A1(_1726_),
    .A2(_1915_),
    .B1_N(_1916_),
    .X(_1999_));
 sky130_fd_sc_hd__nand2_1 _5564_ (.A(net123),
    .B(net148),
    .Y(_2000_));
 sky130_fd_sc_hd__o21ai_1 _5565_ (.A1(net123),
    .A2(net125),
    .B1(net147),
    .Y(_2001_));
 sky130_fd_sc_hd__and3_1 _5566_ (.A(net123),
    .B(net125),
    .C(net147),
    .X(_2002_));
 sky130_fd_sc_hd__nor2_2 _5567_ (.A(_2001_),
    .B(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__xnor2_4 _5568_ (.A(_1823_),
    .B(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__inv_2 _5569_ (.A(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__a32o_1 _5570_ (.A1(net123),
    .A2(net149),
    .A3(_1934_),
    .B1(_1935_),
    .B2(net153),
    .X(_2006_));
 sky130_fd_sc_hd__and2_1 _5571_ (.A(_2004_),
    .B(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__xnor2_1 _5572_ (.A(_2004_),
    .B(_2006_),
    .Y(_2008_));
 sky130_fd_sc_hd__nor2_1 _5573_ (.A(_1999_),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(_1999_),
    .B(_2008_),
    .Y(_2010_));
 sky130_fd_sc_hd__and2b_1 _5575_ (.A_N(_2009_),
    .B(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__xnor2_1 _5576_ (.A(_1998_),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__nor2_1 _5577_ (.A(_1997_),
    .B(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hd__and2_1 _5578_ (.A(_1997_),
    .B(_2012_),
    .X(_2014_));
 sky130_fd_sc_hd__or2_1 _5579_ (.A(_2013_),
    .B(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__a21oi_1 _5580_ (.A1(_1948_),
    .A2(_1951_),
    .B1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__and3_1 _5581_ (.A(_1948_),
    .B(_1951_),
    .C(_2015_),
    .X(_2017_));
 sky130_fd_sc_hd__a211oi_1 _5582_ (.A1(_1924_),
    .A2(_1927_),
    .B1(_2016_),
    .C1(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__o211a_1 _5583_ (.A1(_2016_),
    .A2(_2017_),
    .B1(_1924_),
    .C1(_1927_),
    .X(_2019_));
 sky130_fd_sc_hd__a21o_1 _5584_ (.A1(_1937_),
    .A2(_1946_),
    .B1(_1945_),
    .X(_2020_));
 sky130_fd_sc_hd__nand2_1 _5585_ (.A(net120),
    .B(net150),
    .Y(_2021_));
 sky130_fd_sc_hd__a22o_1 _5586_ (.A1(net115),
    .A2(net155),
    .B1(net152),
    .B2(net117),
    .X(_2022_));
 sky130_fd_sc_hd__and3_1 _5587_ (.A(net115),
    .B(net117),
    .C(net152),
    .X(_2023_));
 sky130_fd_sc_hd__a21bo_1 _5588_ (.A1(net155),
    .A2(_2023_),
    .B1_N(_2022_),
    .X(_2024_));
 sky130_fd_sc_hd__xor2_1 _5589_ (.A(_2021_),
    .B(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__or2_1 _5590_ (.A(_1940_),
    .B(_1943_),
    .X(_2026_));
 sky130_fd_sc_hd__a22oi_1 _5591_ (.A1(\ann.in_ff[2][14] ),
    .A2(net162),
    .B1(net159),
    .B2(net109),
    .Y(_2027_));
 sky130_fd_sc_hd__and4_1 _5592_ (.A(\ann.in_ff[2][14] ),
    .B(net109),
    .C(net162),
    .D(net159),
    .X(_2028_));
 sky130_fd_sc_hd__o2bb2a_1 _5593_ (.A1_N(net112),
    .A2_N(net156),
    .B1(_2027_),
    .B2(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__and4bb_1 _5594_ (.A_N(_2027_),
    .B_N(_2028_),
    .C(net112),
    .D(net156),
    .X(_2030_));
 sky130_fd_sc_hd__nor2_1 _5595_ (.A(_2029_),
    .B(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__nand2_1 _5596_ (.A(_2026_),
    .B(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__xor2_1 _5597_ (.A(_2026_),
    .B(_2031_),
    .X(_2033_));
 sky130_fd_sc_hd__nand2_1 _5598_ (.A(_2025_),
    .B(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__xnor2_1 _5599_ (.A(_2025_),
    .B(_2033_),
    .Y(_2035_));
 sky130_fd_sc_hd__a21o_1 _5600_ (.A1(_1960_),
    .A2(_1962_),
    .B1(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__nand3_1 _5601_ (.A(_1960_),
    .B(_1962_),
    .C(_2035_),
    .Y(_2037_));
 sky130_fd_sc_hd__and3_1 _5602_ (.A(_2020_),
    .B(_2036_),
    .C(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__inv_2 _5603_ (.A(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__a21oi_1 _5604_ (.A1(_2036_),
    .A2(_2037_),
    .B1(_2020_),
    .Y(_2040_));
 sky130_fd_sc_hd__o21ai_1 _5605_ (.A1(_1879_),
    .A2(_1963_),
    .B1(_1878_),
    .Y(_2041_));
 sky130_fd_sc_hd__a31o_1 _5606_ (.A1(\ann.in_ff[2][14] ),
    .A2(net164),
    .A3(_1958_),
    .B1(_1956_),
    .X(_2042_));
 sky130_fd_sc_hd__nand2_2 _5607_ (.A(net105),
    .B(net164),
    .Y(_2043_));
 sky130_fd_sc_hd__xor2_4 _5608_ (.A(_1958_),
    .B(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__nor2_1 _5609_ (.A(_1872_),
    .B(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__xnor2_4 _5610_ (.A(_1872_),
    .B(_2044_),
    .Y(_2046_));
 sky130_fd_sc_hd__and2b_1 _5611_ (.A_N(_2046_),
    .B(_2042_),
    .X(_2047_));
 sky130_fd_sc_hd__xor2_1 _5612_ (.A(_2042_),
    .B(_2046_),
    .X(_2048_));
 sky130_fd_sc_hd__xnor2_1 _5613_ (.A(_1880_),
    .B(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__nand2_1 _5614_ (.A(_2041_),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__or2_1 _5615_ (.A(_2041_),
    .B(_2049_),
    .X(_2051_));
 sky130_fd_sc_hd__nand2_1 _5616_ (.A(_2050_),
    .B(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__or3_1 _5617_ (.A(_2038_),
    .B(_2040_),
    .C(_2052_),
    .X(_2053_));
 sky130_fd_sc_hd__o21ai_1 _5618_ (.A1(_2038_),
    .A2(_2040_),
    .B1(_2052_),
    .Y(_2054_));
 sky130_fd_sc_hd__and2_1 _5619_ (.A(_2053_),
    .B(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__o21ai_2 _5620_ (.A1(_1965_),
    .A2(_1968_),
    .B1(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__or3_1 _5621_ (.A(_1965_),
    .B(_1968_),
    .C(_2055_),
    .X(_2057_));
 sky130_fd_sc_hd__or4bb_4 _5622_ (.A(_2018_),
    .B(_2019_),
    .C_N(_2056_),
    .D_N(_2057_),
    .X(_2058_));
 sky130_fd_sc_hd__a2bb2o_1 _5623_ (.A1_N(_2018_),
    .A2_N(_2019_),
    .B1(_2056_),
    .B2(_2057_),
    .X(_2059_));
 sky130_fd_sc_hd__o211a_1 _5624_ (.A1(_1970_),
    .A2(_1972_),
    .B1(_2058_),
    .C1(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__a211oi_2 _5625_ (.A1(_2058_),
    .A2(_2059_),
    .B1(_1970_),
    .C1(_1972_),
    .Y(_2061_));
 sky130_fd_sc_hd__nor3_1 _5626_ (.A(_1993_),
    .B(_2060_),
    .C(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__or3_1 _5627_ (.A(_1993_),
    .B(_2060_),
    .C(_2061_),
    .X(_2063_));
 sky130_fd_sc_hd__o21ai_1 _5628_ (.A1(_2060_),
    .A2(_2061_),
    .B1(_1993_),
    .Y(_2064_));
 sky130_fd_sc_hd__o211a_1 _5629_ (.A1(_1974_),
    .A2(_1976_),
    .B1(_2063_),
    .C1(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__a211oi_1 _5630_ (.A1(_2063_),
    .A2(_2064_),
    .B1(_1974_),
    .C1(_1976_),
    .Y(_2066_));
 sky130_fd_sc_hd__nor3_1 _5631_ (.A(_1906_),
    .B(_2065_),
    .C(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__o21a_1 _5632_ (.A1(_2065_),
    .A2(_2066_),
    .B1(_1906_),
    .X(_2068_));
 sky130_fd_sc_hd__nor2_1 _5633_ (.A(_2067_),
    .B(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(_1987_),
    .B(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__xnor2_1 _5635_ (.A(_1987_),
    .B(_2069_),
    .Y(_2071_));
 sky130_fd_sc_hd__nand2_1 _5636_ (.A(_1984_),
    .B(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__nor2_1 _5637_ (.A(_1984_),
    .B(_2071_),
    .Y(_2073_));
 sky130_fd_sc_hd__inv_2 _5638_ (.A(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_2072_),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__a2bb2o_1 _5640_ (.A1_N(_1981_),
    .A2_N(_1982_),
    .B1(_1985_),
    .B2(_1903_),
    .X(_2076_));
 sky130_fd_sc_hd__xor2_1 _5641_ (.A(_2075_),
    .B(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__nor2_1 _5642_ (.A(net194),
    .B(_2077_),
    .Y(_0015_));
 sky130_fd_sc_hd__nor2_1 _5643_ (.A(_1276_),
    .B(_1453_),
    .Y(_2078_));
 sky130_fd_sc_hd__nor2_2 _5644_ (.A(_1546_),
    .B(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__a21o_1 _5645_ (.A1(_1725_),
    .A2(_1730_),
    .B1(_1995_),
    .X(_2080_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_2079_),
    .B(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__xor2_2 _5647_ (.A(_2079_),
    .B(_2080_),
    .X(_2082_));
 sky130_fd_sc_hd__nand2b_1 _5648_ (.A_N(_1989_),
    .B(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__xnor2_1 _5649_ (.A(_1989_),
    .B(_2082_),
    .Y(_2084_));
 sky130_fd_sc_hd__or2_1 _5650_ (.A(_2016_),
    .B(_2018_),
    .X(_2085_));
 sky130_fd_sc_hd__nand2_1 _5651_ (.A(_2084_),
    .B(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__xnor2_1 _5652_ (.A(_2084_),
    .B(_2085_),
    .Y(_2087_));
 sky130_fd_sc_hd__a21oi_1 _5653_ (.A1(_1998_),
    .A2(_2011_),
    .B1(_2013_),
    .Y(_2088_));
 sky130_fd_sc_hd__and2b_1 _5654_ (.A_N(_1822_),
    .B(_1827_),
    .X(_2089_));
 sky130_fd_sc_hd__and2b_1 _5655_ (.A_N(_1827_),
    .B(_1822_),
    .X(_2090_));
 sky130_fd_sc_hd__nor2_1 _5656_ (.A(_2089_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__and2_1 _5657_ (.A(_1541_),
    .B(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__nor2_1 _5658_ (.A(_1541_),
    .B(_2091_),
    .Y(_2093_));
 sky130_fd_sc_hd__or2_1 _5659_ (.A(_2092_),
    .B(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__o21ba_2 _5660_ (.A1(_1823_),
    .A2(_2001_),
    .B1_N(_2002_),
    .X(_2095_));
 sky130_fd_sc_hd__nand2_1 _5661_ (.A(net120),
    .B(net148),
    .Y(_2096_));
 sky130_fd_sc_hd__o21ai_1 _5662_ (.A1(net120),
    .A2(net123),
    .B1(net148),
    .Y(_2097_));
 sky130_fd_sc_hd__and3_1 _5663_ (.A(net120),
    .B(net123),
    .C(net148),
    .X(_2098_));
 sky130_fd_sc_hd__nor2_2 _5664_ (.A(_2097_),
    .B(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__xnor2_4 _5665_ (.A(_1914_),
    .B(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__a32o_1 _5666_ (.A1(net120),
    .A2(net150),
    .A3(_2022_),
    .B1(_2023_),
    .B2(net155),
    .X(_2101_));
 sky130_fd_sc_hd__and2_1 _5667_ (.A(_2100_),
    .B(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__xnor2_1 _5668_ (.A(_2100_),
    .B(_2101_),
    .Y(_2103_));
 sky130_fd_sc_hd__nor2_1 _5669_ (.A(_2095_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__xor2_1 _5670_ (.A(_2095_),
    .B(_2103_),
    .X(_2105_));
 sky130_fd_sc_hd__o21ai_1 _5671_ (.A1(_2007_),
    .A2(_2009_),
    .B1(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__or3_1 _5672_ (.A(_2007_),
    .B(_2009_),
    .C(_2105_),
    .X(_2107_));
 sky130_fd_sc_hd__nand2_1 _5673_ (.A(_2106_),
    .B(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__xnor2_1 _5674_ (.A(_2094_),
    .B(_2108_),
    .Y(_2109_));
 sky130_fd_sc_hd__a21oi_1 _5675_ (.A1(_2036_),
    .A2(_2039_),
    .B1(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__and3_1 _5676_ (.A(_2036_),
    .B(_2039_),
    .C(_2109_),
    .X(_2111_));
 sky130_fd_sc_hd__nor3_1 _5677_ (.A(_2088_),
    .B(_2110_),
    .C(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__o21a_1 _5678_ (.A1(_2110_),
    .A2(_2111_),
    .B1(_2088_),
    .X(_2113_));
 sky130_fd_sc_hd__a22o_1 _5679_ (.A1(net111),
    .A2(net155),
    .B1(net152),
    .B2(net114),
    .X(_2114_));
 sky130_fd_sc_hd__and4_1 _5680_ (.A(net111),
    .B(net114),
    .C(net155),
    .D(net152),
    .X(_2115_));
 sky130_fd_sc_hd__inv_2 _5681_ (.A(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__a22oi_1 _5682_ (.A1(net117),
    .A2(net150),
    .B1(_2114_),
    .B2(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__and4b_1 _5683_ (.A_N(_2115_),
    .B(net150),
    .C(net117),
    .D(_2114_),
    .X(_2118_));
 sky130_fd_sc_hd__nor2_1 _5684_ (.A(_2117_),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__or2_1 _5685_ (.A(_2028_),
    .B(_2030_),
    .X(_2120_));
 sky130_fd_sc_hd__nand2_1 _5686_ (.A(net109),
    .B(net156),
    .Y(_2121_));
 sky130_fd_sc_hd__a22oi_1 _5687_ (.A1(net106),
    .A2(net162),
    .B1(net159),
    .B2(net107),
    .Y(_2122_));
 sky130_fd_sc_hd__and4_1 _5688_ (.A(net105),
    .B(net107),
    .C(net162),
    .D(net159),
    .X(_2123_));
 sky130_fd_sc_hd__nor2_1 _5689_ (.A(_2122_),
    .B(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__xnor2_1 _5690_ (.A(_2121_),
    .B(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__and2_1 _5691_ (.A(_2120_),
    .B(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__xor2_1 _5692_ (.A(_2120_),
    .B(_2125_),
    .X(_2127_));
 sky130_fd_sc_hd__xnor2_1 _5693_ (.A(_2119_),
    .B(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__o21bai_2 _5694_ (.A1(_2045_),
    .A2(_2047_),
    .B1_N(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__or3b_1 _5695_ (.A(_2045_),
    .B(_2047_),
    .C_N(_2128_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_1 _5696_ (.A(_2129_),
    .B(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__a21o_1 _5697_ (.A1(_2032_),
    .A2(_2034_),
    .B1(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__nand3_1 _5698_ (.A(_2032_),
    .B(_2034_),
    .C(_2131_),
    .Y(_2133_));
 sky130_fd_sc_hd__o21ai_1 _5699_ (.A1(_1879_),
    .A2(_2048_),
    .B1(_1878_),
    .Y(_2134_));
 sky130_fd_sc_hd__o21ba_1 _5700_ (.A1(_1957_),
    .A2(_2043_),
    .B1_N(_1956_),
    .X(_2135_));
 sky130_fd_sc_hd__xnor2_2 _5701_ (.A(_2046_),
    .B(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__xnor2_1 _5702_ (.A(_1880_),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__and2_1 _5703_ (.A(_2134_),
    .B(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__nor2_1 _5704_ (.A(_2134_),
    .B(_2137_),
    .Y(_2139_));
 sky130_fd_sc_hd__nor2_1 _5705_ (.A(_2138_),
    .B(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__and3_1 _5706_ (.A(_2132_),
    .B(_2133_),
    .C(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__a21oi_1 _5707_ (.A1(_2132_),
    .A2(_2133_),
    .B1(_2140_),
    .Y(_2142_));
 sky130_fd_sc_hd__or2_1 _5708_ (.A(_2141_),
    .B(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__a21oi_2 _5709_ (.A1(_2050_),
    .A2(_2053_),
    .B1(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__and3_1 _5710_ (.A(_2050_),
    .B(_2053_),
    .C(_2143_),
    .X(_2145_));
 sky130_fd_sc_hd__nor4_2 _5711_ (.A(_2112_),
    .B(_2113_),
    .C(_2144_),
    .D(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__o22a_1 _5712_ (.A1(_2112_),
    .A2(_2113_),
    .B1(_2144_),
    .B2(_2145_),
    .X(_2147_));
 sky130_fd_sc_hd__a211oi_2 _5713_ (.A1(_2056_),
    .A2(_2058_),
    .B1(_2146_),
    .C1(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__inv_2 _5714_ (.A(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__o211a_1 _5715_ (.A1(_2146_),
    .A2(_2147_),
    .B1(_2056_),
    .C1(_2058_),
    .X(_2150_));
 sky130_fd_sc_hd__or3_2 _5716_ (.A(_2087_),
    .B(_2148_),
    .C(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__o21ai_2 _5717_ (.A1(_2148_),
    .A2(_2150_),
    .B1(_2087_),
    .Y(_2152_));
 sky130_fd_sc_hd__o211a_1 _5718_ (.A1(_2060_),
    .A2(_2062_),
    .B1(_2151_),
    .C1(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__a211oi_1 _5719_ (.A1(_2151_),
    .A2(_2152_),
    .B1(_2060_),
    .C1(_2062_),
    .Y(_2154_));
 sky130_fd_sc_hd__or3_1 _5720_ (.A(_1992_),
    .B(_2153_),
    .C(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__o21ai_1 _5721_ (.A1(_2153_),
    .A2(_2154_),
    .B1(_1992_),
    .Y(_2156_));
 sky130_fd_sc_hd__o211a_1 _5722_ (.A1(_2065_),
    .A2(_2067_),
    .B1(_2155_),
    .C1(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__a211oi_1 _5723_ (.A1(_2155_),
    .A2(_2156_),
    .B1(_2065_),
    .C1(_2067_),
    .Y(_2158_));
 sky130_fd_sc_hd__nor2_1 _5724_ (.A(_2157_),
    .B(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__and3_1 _5725_ (.A(_1987_),
    .B(_2069_),
    .C(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__xor2_1 _5726_ (.A(_2070_),
    .B(_2159_),
    .X(_2161_));
 sky130_fd_sc_hd__a21oi_2 _5727_ (.A1(_2072_),
    .A2(_2076_),
    .B1(_2073_),
    .Y(_2162_));
 sky130_fd_sc_hd__nor2_1 _5728_ (.A(_2161_),
    .B(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__or2_1 _5729_ (.A(net194),
    .B(_2163_),
    .X(_2164_));
 sky130_fd_sc_hd__a21oi_1 _5730_ (.A1(_2161_),
    .A2(_2162_),
    .B1(_2164_),
    .Y(_0016_));
 sky130_fd_sc_hd__nor2_1 _5731_ (.A(_2160_),
    .B(_2163_),
    .Y(_2165_));
 sky130_fd_sc_hd__nand2b_1 _5732_ (.A_N(_2153_),
    .B(_2155_),
    .Y(_2166_));
 sky130_fd_sc_hd__or2_1 _5733_ (.A(_2110_),
    .B(_2112_),
    .X(_2167_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_1363_),
    .B(_1633_),
    .Y(_2168_));
 sky130_fd_sc_hd__or2_1 _5735_ (.A(_1363_),
    .B(_1633_),
    .X(_2169_));
 sky130_fd_sc_hd__and2_1 _5736_ (.A(_2168_),
    .B(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__o21a_1 _5737_ (.A1(_2089_),
    .A2(_2092_),
    .B1(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__or3_1 _5738_ (.A(_2089_),
    .B(_2092_),
    .C(_2170_),
    .X(_2172_));
 sky130_fd_sc_hd__nand2b_2 _5739_ (.A_N(_2171_),
    .B(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__a21o_1 _5740_ (.A1(_2079_),
    .A2(_2080_),
    .B1(_2078_),
    .X(_2174_));
 sky130_fd_sc_hd__xnor2_2 _5741_ (.A(_2173_),
    .B(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__xnor2_1 _5742_ (.A(_2167_),
    .B(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__and2_1 _5743_ (.A(_2083_),
    .B(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nor2_1 _5744_ (.A(_2083_),
    .B(_2176_),
    .Y(_2178_));
 sky130_fd_sc_hd__o21a_1 _5745_ (.A1(_2094_),
    .A2(_2108_),
    .B1(_2106_),
    .X(_2179_));
 sky130_fd_sc_hd__nand2b_1 _5746_ (.A_N(_1913_),
    .B(_1918_),
    .Y(_2180_));
 sky130_fd_sc_hd__xnor2_2 _5747_ (.A(_1913_),
    .B(_1918_),
    .Y(_2181_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(_1638_),
    .B(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__or2_1 _5749_ (.A(_1638_),
    .B(_2181_),
    .X(_2183_));
 sky130_fd_sc_hd__nand2_1 _5750_ (.A(_2182_),
    .B(_2183_),
    .Y(_2184_));
 sky130_fd_sc_hd__o21ba_1 _5751_ (.A1(_1914_),
    .A2(_2097_),
    .B1_N(_2098_),
    .X(_2185_));
 sky130_fd_sc_hd__and2_1 _5752_ (.A(net117),
    .B(net148),
    .X(_2186_));
 sky130_fd_sc_hd__o21ai_1 _5753_ (.A1(net117),
    .A2(net120),
    .B1(net148),
    .Y(_2187_));
 sky130_fd_sc_hd__and3_1 _5754_ (.A(net117),
    .B(net120),
    .C(net148),
    .X(_2188_));
 sky130_fd_sc_hd__nor2_1 _5755_ (.A(_2187_),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__xnor2_2 _5756_ (.A(_2000_),
    .B(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__or2_1 _5757_ (.A(_2115_),
    .B(_2118_),
    .X(_2191_));
 sky130_fd_sc_hd__and2_1 _5758_ (.A(_2190_),
    .B(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__xnor2_1 _5759_ (.A(_2190_),
    .B(_2191_),
    .Y(_2193_));
 sky130_fd_sc_hd__nor2_1 _5760_ (.A(_2185_),
    .B(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__xor2_1 _5761_ (.A(_2185_),
    .B(_2193_),
    .X(_2195_));
 sky130_fd_sc_hd__o21a_1 _5762_ (.A1(_2102_),
    .A2(_2104_),
    .B1(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__nor3_1 _5763_ (.A(_2102_),
    .B(_2104_),
    .C(_2195_),
    .Y(_2197_));
 sky130_fd_sc_hd__or2_1 _5764_ (.A(_2196_),
    .B(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__nor2_1 _5765_ (.A(_2184_),
    .B(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hd__xnor2_1 _5766_ (.A(_2184_),
    .B(_2198_),
    .Y(_2200_));
 sky130_fd_sc_hd__a21oi_1 _5767_ (.A1(_2129_),
    .A2(_2132_),
    .B1(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__and3_1 _5768_ (.A(_2129_),
    .B(_2132_),
    .C(_2200_),
    .X(_2202_));
 sky130_fd_sc_hd__nor3_1 _5769_ (.A(_2179_),
    .B(_2201_),
    .C(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__o21a_1 _5770_ (.A1(_2201_),
    .A2(_2202_),
    .B1(_2179_),
    .X(_2204_));
 sky130_fd_sc_hd__nor2_1 _5771_ (.A(_2203_),
    .B(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__a31o_1 _5772_ (.A1(_2132_),
    .A2(_2133_),
    .A3(_2140_),
    .B1(_2138_),
    .X(_2206_));
 sky130_fd_sc_hd__a21o_1 _5773_ (.A1(_2119_),
    .A2(_2127_),
    .B1(_2126_),
    .X(_2207_));
 sky130_fd_sc_hd__a22o_1 _5774_ (.A1(net110),
    .A2(net155),
    .B1(net152),
    .B2(net111),
    .X(_2208_));
 sky130_fd_sc_hd__nand4_1 _5775_ (.A(\ann.in_ff[2][13] ),
    .B(net111),
    .C(net155),
    .D(net152),
    .Y(_2209_));
 sky130_fd_sc_hd__a22oi_1 _5776_ (.A1(net114),
    .A2(net150),
    .B1(_2208_),
    .B2(_2209_),
    .Y(_2210_));
 sky130_fd_sc_hd__and4_1 _5777_ (.A(net115),
    .B(net150),
    .C(_2208_),
    .D(_2209_),
    .X(_2211_));
 sky130_fd_sc_hd__nor2_1 _5778_ (.A(_2210_),
    .B(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__a31o_1 _5779_ (.A1(net109),
    .A2(net156),
    .A3(_2124_),
    .B1(_2123_),
    .X(_2213_));
 sky130_fd_sc_hd__nand2_1 _5780_ (.A(net107),
    .B(\ann.weight[11] ),
    .Y(_2214_));
 sky130_fd_sc_hd__o21ai_1 _5781_ (.A1(net162),
    .A2(net159),
    .B1(net105),
    .Y(_2215_));
 sky130_fd_sc_hd__and3_1 _5782_ (.A(net105),
    .B(net162),
    .C(net159),
    .X(_2216_));
 sky130_fd_sc_hd__nor2_1 _5783_ (.A(_2215_),
    .B(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__xnor2_1 _5784_ (.A(_2214_),
    .B(_2217_),
    .Y(_2218_));
 sky130_fd_sc_hd__and2_1 _5785_ (.A(_2213_),
    .B(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__xor2_2 _5786_ (.A(_2213_),
    .B(_2218_),
    .X(_2220_));
 sky130_fd_sc_hd__xnor2_2 _5787_ (.A(_2212_),
    .B(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hd__o21ba_4 _5788_ (.A1(_2046_),
    .A2(_2135_),
    .B1_N(_2045_),
    .X(_2222_));
 sky130_fd_sc_hd__xnor2_1 _5789_ (.A(_2221_),
    .B(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__and2b_1 _5790_ (.A_N(_2223_),
    .B(_2207_),
    .X(_2224_));
 sky130_fd_sc_hd__xnor2_1 _5791_ (.A(_2207_),
    .B(_2223_),
    .Y(_2225_));
 sky130_fd_sc_hd__and2_1 _5792_ (.A(_1879_),
    .B(_2136_),
    .X(_2226_));
 sky130_fd_sc_hd__nor2_4 _5793_ (.A(_1878_),
    .B(_2136_),
    .Y(_2227_));
 sky130_fd_sc_hd__nor2_2 _5794_ (.A(_2226_),
    .B(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__or2_2 _5795_ (.A(_2226_),
    .B(_2227_),
    .X(_2229_));
 sky130_fd_sc_hd__xnor2_1 _5796_ (.A(_2225_),
    .B(_2228_),
    .Y(_2230_));
 sky130_fd_sc_hd__nand2b_1 _5797_ (.A_N(_2230_),
    .B(_2206_),
    .Y(_2231_));
 sky130_fd_sc_hd__nand2b_1 _5798_ (.A_N(_2206_),
    .B(_2230_),
    .Y(_2232_));
 sky130_fd_sc_hd__nand2_1 _5799_ (.A(_2231_),
    .B(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__or3_1 _5800_ (.A(_2203_),
    .B(_2204_),
    .C(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__xnor2_2 _5801_ (.A(_2205_),
    .B(_2233_),
    .Y(_2235_));
 sky130_fd_sc_hd__o21a_1 _5802_ (.A1(_2144_),
    .A2(_2146_),
    .B1(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__nor3_1 _5803_ (.A(_2144_),
    .B(_2146_),
    .C(_2235_),
    .Y(_2237_));
 sky130_fd_sc_hd__nor4_2 _5804_ (.A(_2177_),
    .B(_2178_),
    .C(_2236_),
    .D(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__o22a_1 _5805_ (.A1(_2177_),
    .A2(_2178_),
    .B1(_2236_),
    .B2(_2237_),
    .X(_2239_));
 sky130_fd_sc_hd__a211oi_1 _5806_ (.A1(_2149_),
    .A2(_2151_),
    .B1(_2238_),
    .C1(_2239_),
    .Y(_2240_));
 sky130_fd_sc_hd__o211a_1 _5807_ (.A1(_2238_),
    .A2(_2239_),
    .B1(_2149_),
    .C1(_2151_),
    .X(_2241_));
 sky130_fd_sc_hd__or3_1 _5808_ (.A(_2086_),
    .B(_2240_),
    .C(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__o21ai_1 _5809_ (.A1(_2240_),
    .A2(_2241_),
    .B1(_2086_),
    .Y(_2243_));
 sky130_fd_sc_hd__nand2_2 _5810_ (.A(_2242_),
    .B(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__and2b_1 _5811_ (.A_N(_2244_),
    .B(_2166_),
    .X(_2245_));
 sky130_fd_sc_hd__xnor2_2 _5812_ (.A(_2166_),
    .B(_2244_),
    .Y(_2246_));
 sky130_fd_sc_hd__or2_1 _5813_ (.A(_2157_),
    .B(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__xnor2_1 _5814_ (.A(_2157_),
    .B(_2246_),
    .Y(_2248_));
 sky130_fd_sc_hd__xnor2_1 _5815_ (.A(_2165_),
    .B(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__nor2_1 _5816_ (.A(net194),
    .B(_2249_),
    .Y(_0017_));
 sky130_fd_sc_hd__o21ba_1 _5817_ (.A1(_2086_),
    .A2(_2241_),
    .B1_N(_2240_),
    .X(_2250_));
 sky130_fd_sc_hd__a21oi_2 _5818_ (.A1(_2167_),
    .A2(_2175_),
    .B1(_2178_),
    .Y(_2251_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_1456_),
    .B(_1725_),
    .Y(_2252_));
 sky130_fd_sc_hd__xnor2_1 _5820_ (.A(_1456_),
    .B(_1724_),
    .Y(_2253_));
 sky130_fd_sc_hd__xnor2_1 _5821_ (.A(_1360_),
    .B(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__a21o_1 _5822_ (.A1(_2180_),
    .A2(_2182_),
    .B1(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__nand3_1 _5823_ (.A(_2180_),
    .B(_2182_),
    .C(_2254_),
    .Y(_2256_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_2255_),
    .B(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__xor2_1 _5825_ (.A(_2168_),
    .B(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__o21ai_1 _5826_ (.A1(_2078_),
    .A2(_2171_),
    .B1(_2172_),
    .Y(_2259_));
 sky130_fd_sc_hd__inv_2 _5827_ (.A(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_2258_),
    .B(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__or2_1 _5829_ (.A(_2258_),
    .B(_2260_),
    .X(_2262_));
 sky130_fd_sc_hd__nand2_1 _5830_ (.A(_2261_),
    .B(_2262_),
    .Y(_2263_));
 sky130_fd_sc_hd__nor2_1 _5831_ (.A(_2201_),
    .B(_2203_),
    .Y(_2264_));
 sky130_fd_sc_hd__xnor2_1 _5832_ (.A(_2263_),
    .B(_2264_),
    .Y(_2265_));
 sky130_fd_sc_hd__nor2_1 _5833_ (.A(_2081_),
    .B(_2173_),
    .Y(_2266_));
 sky130_fd_sc_hd__xor2_1 _5834_ (.A(_2265_),
    .B(_2266_),
    .X(_2267_));
 sky130_fd_sc_hd__xnor2_1 _5835_ (.A(_1999_),
    .B(_2004_),
    .Y(_2268_));
 sky130_fd_sc_hd__nand2_1 _5836_ (.A(_1730_),
    .B(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__or2_1 _5837_ (.A(_1730_),
    .B(_2268_),
    .X(_2270_));
 sky130_fd_sc_hd__nand2_1 _5838_ (.A(_2269_),
    .B(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__o21ba_1 _5839_ (.A1(_2000_),
    .A2(_2187_),
    .B1_N(_2188_),
    .X(_2272_));
 sky130_fd_sc_hd__nand2_1 _5840_ (.A(net114),
    .B(net148),
    .Y(_2273_));
 sky130_fd_sc_hd__o21ai_1 _5841_ (.A1(net114),
    .A2(net117),
    .B1(net148),
    .Y(_2274_));
 sky130_fd_sc_hd__and3_1 _5842_ (.A(net114),
    .B(net117),
    .C(net148),
    .X(_2275_));
 sky130_fd_sc_hd__nor2_1 _5843_ (.A(_2274_),
    .B(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__xnor2_2 _5844_ (.A(_2096_),
    .B(_2276_),
    .Y(_2277_));
 sky130_fd_sc_hd__a41o_1 _5845_ (.A1(\ann.in_ff[2][13] ),
    .A2(net111),
    .A3(net155),
    .A4(net152),
    .B1(_2211_),
    .X(_2278_));
 sky130_fd_sc_hd__and2_1 _5846_ (.A(_2277_),
    .B(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__xnor2_1 _5847_ (.A(_2277_),
    .B(_2278_),
    .Y(_2280_));
 sky130_fd_sc_hd__nor2_1 _5848_ (.A(_2272_),
    .B(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__xor2_1 _5849_ (.A(_2272_),
    .B(_2280_),
    .X(_2282_));
 sky130_fd_sc_hd__o21ai_2 _5850_ (.A1(_2192_),
    .A2(_2194_),
    .B1(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__or3_1 _5851_ (.A(_2192_),
    .B(_2194_),
    .C(_2282_),
    .X(_2284_));
 sky130_fd_sc_hd__nand2_1 _5852_ (.A(_2283_),
    .B(_2284_),
    .Y(_2285_));
 sky130_fd_sc_hd__or2_1 _5853_ (.A(_2271_),
    .B(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__xor2_1 _5854_ (.A(_2271_),
    .B(_2285_),
    .X(_2287_));
 sky130_fd_sc_hd__o21bai_2 _5855_ (.A1(_2221_),
    .A2(_2222_),
    .B1_N(_2224_),
    .Y(_2288_));
 sky130_fd_sc_hd__xor2_1 _5856_ (.A(_2287_),
    .B(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__o21a_1 _5857_ (.A1(_2196_),
    .A2(_2199_),
    .B1(_2289_),
    .X(_2290_));
 sky130_fd_sc_hd__nor3_1 _5858_ (.A(_2196_),
    .B(_2199_),
    .C(_2289_),
    .Y(_2291_));
 sky130_fd_sc_hd__a21o_1 _5859_ (.A1(_2225_),
    .A2(_2228_),
    .B1(_2227_),
    .X(_2292_));
 sky130_fd_sc_hd__a21o_1 _5860_ (.A1(_2212_),
    .A2(_2220_),
    .B1(_2219_),
    .X(_2293_));
 sky130_fd_sc_hd__a22oi_1 _5861_ (.A1(net107),
    .A2(net155),
    .B1(net152),
    .B2(net109),
    .Y(_2294_));
 sky130_fd_sc_hd__and4_1 _5862_ (.A(net107),
    .B(net109),
    .C(net155),
    .D(net152),
    .X(_2295_));
 sky130_fd_sc_hd__o2bb2a_1 _5863_ (.A1_N(net112),
    .A2_N(net150),
    .B1(_2294_),
    .B2(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__and4bb_1 _5864_ (.A_N(_2294_),
    .B_N(_2295_),
    .C(net111),
    .D(net150),
    .X(_2297_));
 sky130_fd_sc_hd__nor2_1 _5865_ (.A(_2296_),
    .B(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__a21oi_1 _5866_ (.A1(net107),
    .A2(net157),
    .B1(_2215_),
    .Y(_2299_));
 sky130_fd_sc_hd__or2_1 _5867_ (.A(_2216_),
    .B(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__a21boi_1 _5868_ (.A1(net105),
    .A2(net157),
    .B1_N(_2215_),
    .Y(_2301_));
 sky130_fd_sc_hd__a21oi_1 _5869_ (.A1(net157),
    .A2(_2300_),
    .B1(_2301_),
    .Y(_2302_));
 sky130_fd_sc_hd__xnor2_1 _5870_ (.A(_2298_),
    .B(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__nor2_1 _5871_ (.A(_2222_),
    .B(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__xor2_1 _5872_ (.A(_2222_),
    .B(_2303_),
    .X(_2305_));
 sky130_fd_sc_hd__and2_1 _5873_ (.A(_2293_),
    .B(_2305_),
    .X(_2306_));
 sky130_fd_sc_hd__xnor2_1 _5874_ (.A(_2293_),
    .B(_2305_),
    .Y(_2307_));
 sky130_fd_sc_hd__nor2_1 _5875_ (.A(_2229_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__and2_1 _5876_ (.A(_2229_),
    .B(_2307_),
    .X(_2309_));
 sky130_fd_sc_hd__nor2_1 _5877_ (.A(_2308_),
    .B(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__nand2_1 _5878_ (.A(_2292_),
    .B(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__or2_1 _5879_ (.A(_2292_),
    .B(_2310_),
    .X(_2312_));
 sky130_fd_sc_hd__nand2_1 _5880_ (.A(_2311_),
    .B(_2312_),
    .Y(_2313_));
 sky130_fd_sc_hd__nor3_1 _5881_ (.A(_2290_),
    .B(_2291_),
    .C(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__or3_1 _5882_ (.A(_2290_),
    .B(_2291_),
    .C(_2313_),
    .X(_2315_));
 sky130_fd_sc_hd__o21a_1 _5883_ (.A1(_2290_),
    .A2(_2291_),
    .B1(_2313_),
    .X(_2316_));
 sky130_fd_sc_hd__a211oi_2 _5884_ (.A1(_2231_),
    .A2(_2234_),
    .B1(_2314_),
    .C1(_2316_),
    .Y(_2317_));
 sky130_fd_sc_hd__o211a_1 _5885_ (.A1(_2314_),
    .A2(_2316_),
    .B1(_2231_),
    .C1(_2234_),
    .X(_2318_));
 sky130_fd_sc_hd__or3_1 _5886_ (.A(_2267_),
    .B(_2317_),
    .C(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__o21ai_1 _5887_ (.A1(_2317_),
    .A2(_2318_),
    .B1(_2267_),
    .Y(_2320_));
 sky130_fd_sc_hd__o211a_1 _5888_ (.A1(_2236_),
    .A2(_2238_),
    .B1(_2319_),
    .C1(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__a211o_1 _5889_ (.A1(_2319_),
    .A2(_2320_),
    .B1(_2236_),
    .C1(_2238_),
    .X(_2322_));
 sky130_fd_sc_hd__and2b_1 _5890_ (.A_N(_2321_),
    .B(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__or3b_1 _5891_ (.A(_2251_),
    .B(_2321_),
    .C_N(_2322_),
    .X(_2324_));
 sky130_fd_sc_hd__xnor2_2 _5892_ (.A(_2251_),
    .B(_2323_),
    .Y(_2325_));
 sky130_fd_sc_hd__and2b_1 _5893_ (.A_N(_2250_),
    .B(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__xnor2_2 _5894_ (.A(_2250_),
    .B(_2325_),
    .Y(_2327_));
 sky130_fd_sc_hd__and2_1 _5895_ (.A(_2245_),
    .B(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__xor2_2 _5896_ (.A(_2245_),
    .B(_2327_),
    .X(_2329_));
 sky130_fd_sc_hd__o21a_1 _5897_ (.A1(_2157_),
    .A2(_2160_),
    .B1(_2246_),
    .X(_2330_));
 sky130_fd_sc_hd__a21o_1 _5898_ (.A1(_2163_),
    .A2(_2247_),
    .B1(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__or2_1 _5899_ (.A(_2329_),
    .B(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__nand2_1 _5900_ (.A(_2329_),
    .B(_2331_),
    .Y(_2333_));
 sky130_fd_sc_hd__and3_1 _5901_ (.A(net198),
    .B(_2332_),
    .C(_2333_),
    .X(_0018_));
 sky130_fd_sc_hd__a21o_1 _5902_ (.A1(_2329_),
    .A2(_2331_),
    .B1(_2328_),
    .X(_2334_));
 sky130_fd_sc_hd__and2b_1 _5903_ (.A_N(_2321_),
    .B(_2324_),
    .X(_2335_));
 sky130_fd_sc_hd__o32a_1 _5904_ (.A1(_2081_),
    .A2(_2173_),
    .A3(_2265_),
    .B1(_2264_),
    .B2(_2263_),
    .X(_2336_));
 sky130_fd_sc_hd__and2b_1 _5905_ (.A_N(_2317_),
    .B(_2319_),
    .X(_2337_));
 sky130_fd_sc_hd__o21ai_2 _5906_ (.A1(_2168_),
    .A2(_2257_),
    .B1(_2255_),
    .Y(_2338_));
 sky130_fd_sc_hd__a21bo_1 _5907_ (.A1(_1360_),
    .A2(_2253_),
    .B1_N(_2252_),
    .X(_2339_));
 sky130_fd_sc_hd__nor2_1 _5908_ (.A(_1542_),
    .B(_1822_),
    .Y(_2340_));
 sky130_fd_sc_hd__and2_1 _5909_ (.A(_1542_),
    .B(_1822_),
    .X(_2341_));
 sky130_fd_sc_hd__nor2_1 _5910_ (.A(_2340_),
    .B(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__xor2_1 _5911_ (.A(_1547_),
    .B(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__o21a_1 _5912_ (.A1(_1999_),
    .A2(_2005_),
    .B1(_2269_),
    .X(_2344_));
 sky130_fd_sc_hd__and2b_1 _5913_ (.A_N(_2344_),
    .B(_2343_),
    .X(_2345_));
 sky130_fd_sc_hd__xor2_1 _5914_ (.A(_2343_),
    .B(_2344_),
    .X(_2346_));
 sky130_fd_sc_hd__and2b_1 _5915_ (.A_N(_2346_),
    .B(_2339_),
    .X(_2347_));
 sky130_fd_sc_hd__xnor2_1 _5916_ (.A(_2339_),
    .B(_2346_),
    .Y(_2348_));
 sky130_fd_sc_hd__xnor2_1 _5917_ (.A(_2338_),
    .B(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__or2_1 _5918_ (.A(_1276_),
    .B(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_1276_),
    .B(_2349_),
    .Y(_2351_));
 sky130_fd_sc_hd__and2_1 _5920_ (.A(_2350_),
    .B(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__a21oi_1 _5921_ (.A1(_2287_),
    .A2(_2288_),
    .B1(_2290_),
    .Y(_2353_));
 sky130_fd_sc_hd__nand2b_1 _5922_ (.A_N(_2353_),
    .B(_2352_),
    .Y(_2354_));
 sky130_fd_sc_hd__xnor2_1 _5923_ (.A(_2352_),
    .B(_2353_),
    .Y(_2355_));
 sky130_fd_sc_hd__nand2b_1 _5924_ (.A_N(_2261_),
    .B(_2355_),
    .Y(_2356_));
 sky130_fd_sc_hd__xnor2_1 _5925_ (.A(_2261_),
    .B(_2355_),
    .Y(_2357_));
 sky130_fd_sc_hd__and2b_1 _5926_ (.A_N(_2095_),
    .B(_2100_),
    .X(_2358_));
 sky130_fd_sc_hd__and2b_1 _5927_ (.A_N(_2100_),
    .B(_2095_),
    .X(_2359_));
 sky130_fd_sc_hd__nor2_1 _5928_ (.A(_2358_),
    .B(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__xnor2_2 _5929_ (.A(_1827_),
    .B(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__o21ba_1 _5930_ (.A1(_2096_),
    .A2(_2274_),
    .B1_N(_2275_),
    .X(_2362_));
 sky130_fd_sc_hd__nand2_1 _5931_ (.A(net111),
    .B(net148),
    .Y(_2363_));
 sky130_fd_sc_hd__o21ai_1 _5932_ (.A1(net111),
    .A2(net114),
    .B1(net148),
    .Y(_2364_));
 sky130_fd_sc_hd__and3_1 _5933_ (.A(net111),
    .B(net114),
    .C(\ann.weight[15] ),
    .X(_2365_));
 sky130_fd_sc_hd__nor2_1 _5934_ (.A(_2364_),
    .B(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__xor2_2 _5935_ (.A(_2186_),
    .B(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__or2_1 _5936_ (.A(_2295_),
    .B(_2297_),
    .X(_2368_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(_2367_),
    .B(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__xnor2_1 _5938_ (.A(_2367_),
    .B(_2368_),
    .Y(_2370_));
 sky130_fd_sc_hd__xor2_1 _5939_ (.A(_2362_),
    .B(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__o21ai_1 _5940_ (.A1(_2279_),
    .A2(_2281_),
    .B1(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__or3_1 _5941_ (.A(_2279_),
    .B(_2281_),
    .C(_2371_),
    .X(_2373_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_2372_),
    .B(_2373_),
    .Y(_2374_));
 sky130_fd_sc_hd__or2_1 _5943_ (.A(_2361_),
    .B(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__xor2_1 _5944_ (.A(_2361_),
    .B(_2374_),
    .X(_2376_));
 sky130_fd_sc_hd__o21ai_1 _5945_ (.A1(_2304_),
    .A2(_2306_),
    .B1(_2376_),
    .Y(_2377_));
 sky130_fd_sc_hd__or3_1 _5946_ (.A(_2304_),
    .B(_2306_),
    .C(_2376_),
    .X(_2378_));
 sky130_fd_sc_hd__nand2_1 _5947_ (.A(_2377_),
    .B(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__a21o_1 _5948_ (.A1(_2283_),
    .A2(_2286_),
    .B1(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__nand3_1 _5949_ (.A(_2283_),
    .B(_2286_),
    .C(_2379_),
    .Y(_2381_));
 sky130_fd_sc_hd__and2_1 _5950_ (.A(net157),
    .B(_2216_),
    .X(_2382_));
 sky130_fd_sc_hd__nand2_1 _5951_ (.A(net157),
    .B(_2216_),
    .Y(_2383_));
 sky130_fd_sc_hd__a21o_1 _5952_ (.A1(_2298_),
    .A2(_2302_),
    .B1(_2382_),
    .X(_2384_));
 sky130_fd_sc_hd__a22oi_1 _5953_ (.A1(net105),
    .A2(net155),
    .B1(net152),
    .B2(net107),
    .Y(_2385_));
 sky130_fd_sc_hd__and4_1 _5954_ (.A(net105),
    .B(net107),
    .C(net155),
    .D(net152),
    .X(_2386_));
 sky130_fd_sc_hd__nor2_1 _5955_ (.A(_2385_),
    .B(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__a21oi_1 _5956_ (.A1(net109),
    .A2(net150),
    .B1(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__and3_1 _5957_ (.A(net109),
    .B(net150),
    .C(_2387_),
    .X(_2389_));
 sky130_fd_sc_hd__or2_1 _5958_ (.A(_2388_),
    .B(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__or2_4 _5959_ (.A(_2301_),
    .B(_2382_),
    .X(_2391_));
 sky130_fd_sc_hd__xor2_1 _5960_ (.A(_2390_),
    .B(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__nand2b_1 _5961_ (.A_N(_2222_),
    .B(_2392_),
    .Y(_2393_));
 sky130_fd_sc_hd__xor2_1 _5962_ (.A(_2222_),
    .B(_2392_),
    .X(_2394_));
 sky130_fd_sc_hd__nand2b_1 _5963_ (.A_N(_2394_),
    .B(_2384_),
    .Y(_2395_));
 sky130_fd_sc_hd__xor2_1 _5964_ (.A(_2384_),
    .B(_2394_),
    .X(_2396_));
 sky130_fd_sc_hd__nor2_1 _5965_ (.A(_2229_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__and2_1 _5966_ (.A(_2229_),
    .B(_2396_),
    .X(_2398_));
 sky130_fd_sc_hd__nor2_1 _5967_ (.A(_2397_),
    .B(_2398_),
    .Y(_2399_));
 sky130_fd_sc_hd__o21a_1 _5968_ (.A1(_2227_),
    .A2(_2308_),
    .B1(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__nor3_1 _5969_ (.A(_2227_),
    .B(_2308_),
    .C(_2399_),
    .Y(_2401_));
 sky130_fd_sc_hd__nor2_1 _5970_ (.A(_2400_),
    .B(_2401_),
    .Y(_2402_));
 sky130_fd_sc_hd__and3_1 _5971_ (.A(_2380_),
    .B(_2381_),
    .C(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__a21oi_1 _5972_ (.A1(_2380_),
    .A2(_2381_),
    .B1(_2402_),
    .Y(_2404_));
 sky130_fd_sc_hd__a211o_1 _5973_ (.A1(_2311_),
    .A2(_2315_),
    .B1(_2403_),
    .C1(_2404_),
    .X(_2405_));
 sky130_fd_sc_hd__o211ai_1 _5974_ (.A1(_2403_),
    .A2(_2404_),
    .B1(_2311_),
    .C1(_2315_),
    .Y(_2406_));
 sky130_fd_sc_hd__nand3_1 _5975_ (.A(_2357_),
    .B(_2405_),
    .C(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__a21o_1 _5976_ (.A1(_2405_),
    .A2(_2406_),
    .B1(_2357_),
    .X(_2408_));
 sky130_fd_sc_hd__nand2_2 _5977_ (.A(_2407_),
    .B(_2408_),
    .Y(_2409_));
 sky130_fd_sc_hd__xor2_2 _5978_ (.A(_2337_),
    .B(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__and2b_1 _5979_ (.A_N(_2336_),
    .B(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__xnor2_2 _5980_ (.A(_2336_),
    .B(_2410_),
    .Y(_2412_));
 sky130_fd_sc_hd__and2b_1 _5981_ (.A_N(_2335_),
    .B(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__xnor2_2 _5982_ (.A(_2335_),
    .B(_2412_),
    .Y(_2414_));
 sky130_fd_sc_hd__xor2_2 _5983_ (.A(_2326_),
    .B(_2414_),
    .X(_2415_));
 sky130_fd_sc_hd__xnor2_1 _5984_ (.A(_2334_),
    .B(_2415_),
    .Y(_2416_));
 sky130_fd_sc_hd__nor2_1 _5985_ (.A(net194),
    .B(_2416_),
    .Y(_0019_));
 sky130_fd_sc_hd__and4bb_1 _5986_ (.A_N(_2161_),
    .B_N(_2248_),
    .C(_2329_),
    .D(_2415_),
    .X(_2417_));
 sky130_fd_sc_hd__inv_2 _5987_ (.A(_2417_),
    .Y(_2418_));
 sky130_fd_sc_hd__o21a_1 _5988_ (.A1(_2326_),
    .A2(_2328_),
    .B1(_2414_),
    .X(_2419_));
 sky130_fd_sc_hd__a31o_1 _5989_ (.A1(_2329_),
    .A2(_2330_),
    .A3(_2415_),
    .B1(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__o21bai_2 _5990_ (.A1(_2162_),
    .A2(_2418_),
    .B1_N(_2420_),
    .Y(_2421_));
 sky130_fd_sc_hd__o21ba_1 _5991_ (.A1(_2337_),
    .A2(_2409_),
    .B1_N(_2411_),
    .X(_2422_));
 sky130_fd_sc_hd__nand2_1 _5992_ (.A(_2405_),
    .B(_2407_),
    .Y(_2423_));
 sky130_fd_sc_hd__a21bo_1 _5993_ (.A1(_2338_),
    .A2(_2348_),
    .B1_N(_2350_),
    .X(_2424_));
 sky130_fd_sc_hd__a21oi_1 _5994_ (.A1(_1547_),
    .A2(_2342_),
    .B1(_2340_),
    .Y(_2425_));
 sky130_fd_sc_hd__and2b_1 _5995_ (.A_N(_1913_),
    .B(_1638_),
    .X(_2426_));
 sky130_fd_sc_hd__and2b_1 _5996_ (.A_N(_1638_),
    .B(_1913_),
    .X(_2427_));
 sky130_fd_sc_hd__nor2_1 _5997_ (.A(_2426_),
    .B(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__xnor2_2 _5998_ (.A(_1632_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__a21oi_1 _5999_ (.A1(_1827_),
    .A2(_2360_),
    .B1(_2358_),
    .Y(_2430_));
 sky130_fd_sc_hd__and2b_1 _6000_ (.A_N(_2430_),
    .B(_2429_),
    .X(_2431_));
 sky130_fd_sc_hd__xnor2_1 _6001_ (.A(_2429_),
    .B(_2430_),
    .Y(_2432_));
 sky130_fd_sc_hd__and2b_1 _6002_ (.A_N(_2425_),
    .B(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__xnor2_1 _6003_ (.A(_2425_),
    .B(_2432_),
    .Y(_2434_));
 sky130_fd_sc_hd__o21a_1 _6004_ (.A1(_2345_),
    .A2(_2347_),
    .B1(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__nor3_1 _6005_ (.A(_2345_),
    .B(_2347_),
    .C(_2434_),
    .Y(_2436_));
 sky130_fd_sc_hd__nor2_1 _6006_ (.A(_2435_),
    .B(_2436_),
    .Y(_2437_));
 sky130_fd_sc_hd__xnor2_1 _6007_ (.A(_1363_),
    .B(_2437_),
    .Y(_2438_));
 sky130_fd_sc_hd__a21oi_1 _6008_ (.A1(_2377_),
    .A2(_2380_),
    .B1(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__and3_1 _6009_ (.A(_2377_),
    .B(_2380_),
    .C(_2438_),
    .X(_2440_));
 sky130_fd_sc_hd__nor2_1 _6010_ (.A(_2439_),
    .B(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__xor2_1 _6011_ (.A(_2424_),
    .B(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__and2b_1 _6012_ (.A_N(_2185_),
    .B(_2190_),
    .X(_2443_));
 sky130_fd_sc_hd__and2b_1 _6013_ (.A_N(_2190_),
    .B(_2185_),
    .X(_2444_));
 sky130_fd_sc_hd__nor2_1 _6014_ (.A(_2443_),
    .B(_2444_),
    .Y(_2445_));
 sky130_fd_sc_hd__and2_1 _6015_ (.A(_1918_),
    .B(_2445_),
    .X(_2446_));
 sky130_fd_sc_hd__nor2_1 _6016_ (.A(_1918_),
    .B(_2445_),
    .Y(_2447_));
 sky130_fd_sc_hd__or2_1 _6017_ (.A(_2446_),
    .B(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__o21ai_2 _6018_ (.A1(_2362_),
    .A2(_2370_),
    .B1(_2369_),
    .Y(_2449_));
 sky130_fd_sc_hd__a21o_1 _6019_ (.A1(_2186_),
    .A2(_2366_),
    .B1(_2365_),
    .X(_2450_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(net109),
    .B(\ann.weight[15] ),
    .Y(_2451_));
 sky130_fd_sc_hd__and2_1 _6021_ (.A(_2363_),
    .B(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__nor2_1 _6022_ (.A(_2363_),
    .B(_2451_),
    .Y(_2453_));
 sky130_fd_sc_hd__nor2_1 _6023_ (.A(_2452_),
    .B(_2453_),
    .Y(_2454_));
 sky130_fd_sc_hd__xnor2_2 _6024_ (.A(_2273_),
    .B(_2454_),
    .Y(_2455_));
 sky130_fd_sc_hd__nor2_1 _6025_ (.A(_2386_),
    .B(_2389_),
    .Y(_2456_));
 sky130_fd_sc_hd__and2b_1 _6026_ (.A_N(_2456_),
    .B(_2455_),
    .X(_2457_));
 sky130_fd_sc_hd__xnor2_1 _6027_ (.A(_2455_),
    .B(_2456_),
    .Y(_2458_));
 sky130_fd_sc_hd__xor2_1 _6028_ (.A(_2450_),
    .B(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__nand2_1 _6029_ (.A(_2449_),
    .B(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__xnor2_1 _6030_ (.A(_2449_),
    .B(_2459_),
    .Y(_2461_));
 sky130_fd_sc_hd__or2_1 _6031_ (.A(_2448_),
    .B(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__xnor2_1 _6032_ (.A(_2448_),
    .B(_2461_),
    .Y(_2463_));
 sky130_fd_sc_hd__a21oi_1 _6033_ (.A1(_2393_),
    .A2(_2395_),
    .B1(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__and3_1 _6034_ (.A(_2393_),
    .B(_2395_),
    .C(_2463_),
    .X(_2465_));
 sky130_fd_sc_hd__a211oi_1 _6035_ (.A1(_2372_),
    .A2(_2375_),
    .B1(_2464_),
    .C1(_2465_),
    .Y(_2466_));
 sky130_fd_sc_hd__o211ai_1 _6036_ (.A1(_2464_),
    .A2(_2465_),
    .B1(_2372_),
    .C1(_2375_),
    .Y(_2467_));
 sky130_fd_sc_hd__and2b_1 _6037_ (.A_N(_2466_),
    .B(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__o21ai_2 _6038_ (.A1(_2390_),
    .A2(_2391_),
    .B1(_2383_),
    .Y(_2469_));
 sky130_fd_sc_hd__nand2_1 _6039_ (.A(net107),
    .B(net150),
    .Y(_2470_));
 sky130_fd_sc_hd__and3_1 _6040_ (.A(net105),
    .B(net155),
    .C(\ann.weight[13] ),
    .X(_2471_));
 sky130_fd_sc_hd__o21ai_1 _6041_ (.A1(net155),
    .A2(\ann.weight[13] ),
    .B1(net105),
    .Y(_2472_));
 sky130_fd_sc_hd__nor2_1 _6042_ (.A(_2471_),
    .B(_2472_),
    .Y(_2473_));
 sky130_fd_sc_hd__xnor2_1 _6043_ (.A(_2470_),
    .B(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__and2b_1 _6044_ (.A_N(_2391_),
    .B(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__xnor2_1 _6045_ (.A(_2391_),
    .B(_2474_),
    .Y(_2476_));
 sky130_fd_sc_hd__nand2b_1 _6046_ (.A_N(_2222_),
    .B(_2476_),
    .Y(_2477_));
 sky130_fd_sc_hd__xnor2_1 _6047_ (.A(_2222_),
    .B(_2476_),
    .Y(_2478_));
 sky130_fd_sc_hd__xnor2_1 _6048_ (.A(_2469_),
    .B(_2478_),
    .Y(_2479_));
 sky130_fd_sc_hd__nor2_1 _6049_ (.A(_2229_),
    .B(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__and2_1 _6050_ (.A(_2229_),
    .B(_2479_),
    .X(_2481_));
 sky130_fd_sc_hd__nor2_1 _6051_ (.A(_2480_),
    .B(_2481_),
    .Y(_2482_));
 sky130_fd_sc_hd__o21a_1 _6052_ (.A1(_2227_),
    .A2(_2397_),
    .B1(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__nor3_1 _6053_ (.A(_2227_),
    .B(_2397_),
    .C(_2482_),
    .Y(_2484_));
 sky130_fd_sc_hd__nor2_1 _6054_ (.A(_2483_),
    .B(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__and2_1 _6055_ (.A(_2468_),
    .B(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__nor2_1 _6056_ (.A(_2468_),
    .B(_2485_),
    .Y(_2487_));
 sky130_fd_sc_hd__nor2_1 _6057_ (.A(_2486_),
    .B(_2487_),
    .Y(_2488_));
 sky130_fd_sc_hd__o21ai_1 _6058_ (.A1(_2400_),
    .A2(_2403_),
    .B1(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__or3_1 _6059_ (.A(_2400_),
    .B(_2403_),
    .C(_2488_),
    .X(_2490_));
 sky130_fd_sc_hd__nand3_1 _6060_ (.A(_2442_),
    .B(_2489_),
    .C(_2490_),
    .Y(_2491_));
 sky130_fd_sc_hd__a21o_1 _6061_ (.A1(_2489_),
    .A2(_2490_),
    .B1(_2442_),
    .X(_2492_));
 sky130_fd_sc_hd__and3_1 _6062_ (.A(_2423_),
    .B(_2491_),
    .C(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__a21oi_1 _6063_ (.A1(_2491_),
    .A2(_2492_),
    .B1(_2423_),
    .Y(_2494_));
 sky130_fd_sc_hd__a211oi_1 _6064_ (.A1(_2354_),
    .A2(_2356_),
    .B1(_2493_),
    .C1(_2494_),
    .Y(_2495_));
 sky130_fd_sc_hd__o211ai_1 _6065_ (.A1(_2493_),
    .A2(_2494_),
    .B1(_2354_),
    .C1(_2356_),
    .Y(_2496_));
 sky130_fd_sc_hd__and2b_2 _6066_ (.A_N(_2495_),
    .B(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__and2b_1 _6067_ (.A_N(_2422_),
    .B(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__xnor2_1 _6068_ (.A(_2422_),
    .B(_2497_),
    .Y(_2499_));
 sky130_fd_sc_hd__and2_1 _6069_ (.A(_2413_),
    .B(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__nor2_1 _6070_ (.A(_2413_),
    .B(_2499_),
    .Y(_2501_));
 sky130_fd_sc_hd__nor2_1 _6071_ (.A(_2500_),
    .B(_2501_),
    .Y(_2502_));
 sky130_fd_sc_hd__a21oi_1 _6072_ (.A1(_2421_),
    .A2(_2502_),
    .B1(net195),
    .Y(_2503_));
 sky130_fd_sc_hd__o21a_1 _6073_ (.A1(_2421_),
    .A2(_2502_),
    .B1(_2503_),
    .X(_0020_));
 sky130_fd_sc_hd__a21o_1 _6074_ (.A1(_2421_),
    .A2(_2502_),
    .B1(_2500_),
    .X(_2504_));
 sky130_fd_sc_hd__or2_2 _6075_ (.A(_2493_),
    .B(_2495_),
    .X(_2505_));
 sky130_fd_sc_hd__a21oi_1 _6076_ (.A1(_2424_),
    .A2(_2441_),
    .B1(_2439_),
    .Y(_2506_));
 sky130_fd_sc_hd__nand2_1 _6077_ (.A(_2489_),
    .B(_2491_),
    .Y(_2507_));
 sky130_fd_sc_hd__a21oi_2 _6078_ (.A1(_1363_),
    .A2(_2437_),
    .B1(_2435_),
    .Y(_2508_));
 sky130_fd_sc_hd__or2_1 _6079_ (.A(_2431_),
    .B(_2433_),
    .X(_2509_));
 sky130_fd_sc_hd__a21oi_2 _6080_ (.A1(_1633_),
    .A2(_2428_),
    .B1(_2426_),
    .Y(_2510_));
 sky130_fd_sc_hd__nand2b_1 _6081_ (.A_N(_1999_),
    .B(_1730_),
    .Y(_2511_));
 sky130_fd_sc_hd__xnor2_1 _6082_ (.A(_1730_),
    .B(_1999_),
    .Y(_2512_));
 sky130_fd_sc_hd__xnor2_1 _6083_ (.A(_1724_),
    .B(_2512_),
    .Y(_2513_));
 sky130_fd_sc_hd__o21a_1 _6084_ (.A1(_2443_),
    .A2(_2446_),
    .B1(_2513_),
    .X(_2514_));
 sky130_fd_sc_hd__nor3_1 _6085_ (.A(_2443_),
    .B(_2446_),
    .C(_2513_),
    .Y(_2515_));
 sky130_fd_sc_hd__nor2_1 _6086_ (.A(_2514_),
    .B(_2515_),
    .Y(_2516_));
 sky130_fd_sc_hd__and2b_1 _6087_ (.A_N(_2510_),
    .B(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__xnor2_1 _6088_ (.A(_2510_),
    .B(_2516_),
    .Y(_2518_));
 sky130_fd_sc_hd__xnor2_1 _6089_ (.A(_2509_),
    .B(_2518_),
    .Y(_2519_));
 sky130_fd_sc_hd__nor2_1 _6090_ (.A(_1723_),
    .B(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__and2_1 _6091_ (.A(_1723_),
    .B(_2519_),
    .X(_2521_));
 sky130_fd_sc_hd__nor2_1 _6092_ (.A(_2520_),
    .B(_2521_),
    .Y(_2522_));
 sky130_fd_sc_hd__or2_1 _6093_ (.A(_2464_),
    .B(_2466_),
    .X(_2523_));
 sky130_fd_sc_hd__xnor2_1 _6094_ (.A(_2522_),
    .B(_2523_),
    .Y(_2524_));
 sky130_fd_sc_hd__nor2_1 _6095_ (.A(_2508_),
    .B(_2524_),
    .Y(_2525_));
 sky130_fd_sc_hd__and2_1 _6096_ (.A(_2508_),
    .B(_2524_),
    .X(_2526_));
 sky130_fd_sc_hd__and2b_1 _6097_ (.A_N(_2272_),
    .B(_2277_),
    .X(_2527_));
 sky130_fd_sc_hd__and2b_1 _6098_ (.A_N(_2277_),
    .B(_2272_),
    .X(_2528_));
 sky130_fd_sc_hd__or2_1 _6099_ (.A(_2527_),
    .B(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__nor2_1 _6100_ (.A(_2005_),
    .B(_2529_),
    .Y(_2530_));
 sky130_fd_sc_hd__and2_1 _6101_ (.A(_2005_),
    .B(_2529_),
    .X(_2531_));
 sky130_fd_sc_hd__or2_1 _6102_ (.A(_2530_),
    .B(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__a21o_1 _6103_ (.A1(_2450_),
    .A2(_2458_),
    .B1(_2457_),
    .X(_2533_));
 sky130_fd_sc_hd__a31o_1 _6104_ (.A1(net114),
    .A2(net148),
    .A3(_2454_),
    .B1(_2453_),
    .X(_2534_));
 sky130_fd_sc_hd__and3_1 _6105_ (.A(net107),
    .B(net109),
    .C(\ann.weight[15] ),
    .X(_2535_));
 sky130_fd_sc_hd__or2_1 _6106_ (.A(net107),
    .B(net109),
    .X(_2536_));
 sky130_fd_sc_hd__and3b_1 _6107_ (.A_N(_2535_),
    .B(_2536_),
    .C(\ann.weight[15] ),
    .X(_2537_));
 sky130_fd_sc_hd__mux2_1 _6108_ (.A0(_2363_),
    .A1(net111),
    .S(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__a31o_1 _6109_ (.A1(net107),
    .A2(net150),
    .A3(_2473_),
    .B1(_2471_),
    .X(_2539_));
 sky130_fd_sc_hd__nand2b_1 _6110_ (.A_N(_2538_),
    .B(_2539_),
    .Y(_2540_));
 sky130_fd_sc_hd__xor2_1 _6111_ (.A(_2538_),
    .B(_2539_),
    .X(_2541_));
 sky130_fd_sc_hd__nand2b_1 _6112_ (.A_N(_2541_),
    .B(_2534_),
    .Y(_2542_));
 sky130_fd_sc_hd__xnor2_1 _6113_ (.A(_2534_),
    .B(_2541_),
    .Y(_2543_));
 sky130_fd_sc_hd__nand2_1 _6114_ (.A(_2533_),
    .B(_2543_),
    .Y(_2544_));
 sky130_fd_sc_hd__xnor2_1 _6115_ (.A(_2533_),
    .B(_2543_),
    .Y(_2545_));
 sky130_fd_sc_hd__or2_2 _6116_ (.A(_2532_),
    .B(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__nand2_1 _6117_ (.A(_2532_),
    .B(_2545_),
    .Y(_2547_));
 sky130_fd_sc_hd__a21bo_1 _6118_ (.A1(_2469_),
    .A2(_2478_),
    .B1_N(_2477_),
    .X(_2548_));
 sky130_fd_sc_hd__and3_1 _6119_ (.A(_2546_),
    .B(_2547_),
    .C(_2548_),
    .X(_2549_));
 sky130_fd_sc_hd__a21oi_1 _6120_ (.A1(_2546_),
    .A2(_2547_),
    .B1(_2548_),
    .Y(_2550_));
 sky130_fd_sc_hd__or2_1 _6121_ (.A(_2549_),
    .B(_2550_),
    .X(_2551_));
 sky130_fd_sc_hd__a21oi_2 _6122_ (.A1(_2460_),
    .A2(_2462_),
    .B1(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__and3_1 _6123_ (.A(_2460_),
    .B(_2462_),
    .C(_2551_),
    .X(_2553_));
 sky130_fd_sc_hd__a21oi_1 _6124_ (.A1(net105),
    .A2(net150),
    .B1(_2473_),
    .Y(_2554_));
 sky130_fd_sc_hd__and2_1 _6125_ (.A(net150),
    .B(_2473_),
    .X(_2555_));
 sky130_fd_sc_hd__or2_1 _6126_ (.A(_2554_),
    .B(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__xor2_2 _6127_ (.A(_2391_),
    .B(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__nand2b_1 _6128_ (.A_N(_2222_),
    .B(_2557_),
    .Y(_2558_));
 sky130_fd_sc_hd__xnor2_2 _6129_ (.A(_2222_),
    .B(_2557_),
    .Y(_2559_));
 sky130_fd_sc_hd__o21ai_1 _6130_ (.A1(_2382_),
    .A2(_2475_),
    .B1(_2559_),
    .Y(_2560_));
 sky130_fd_sc_hd__or3_1 _6131_ (.A(_2382_),
    .B(_2475_),
    .C(_2559_),
    .X(_2561_));
 sky130_fd_sc_hd__nand2_1 _6132_ (.A(_2560_),
    .B(_2561_),
    .Y(_2562_));
 sky130_fd_sc_hd__nor2_1 _6133_ (.A(_2229_),
    .B(_2562_),
    .Y(_2563_));
 sky130_fd_sc_hd__and2_1 _6134_ (.A(_2229_),
    .B(_2562_),
    .X(_2564_));
 sky130_fd_sc_hd__nor2_1 _6135_ (.A(_2563_),
    .B(_2564_),
    .Y(_2565_));
 sky130_fd_sc_hd__o21a_1 _6136_ (.A1(_2227_),
    .A2(_2480_),
    .B1(_2565_),
    .X(_2566_));
 sky130_fd_sc_hd__nor3_1 _6137_ (.A(_2227_),
    .B(_2480_),
    .C(_2565_),
    .Y(_2567_));
 sky130_fd_sc_hd__or2_1 _6138_ (.A(_2566_),
    .B(_2567_),
    .X(_2568_));
 sky130_fd_sc_hd__nor3_1 _6139_ (.A(_2552_),
    .B(_2553_),
    .C(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__o21a_1 _6140_ (.A1(_2552_),
    .A2(_2553_),
    .B1(_2568_),
    .X(_2570_));
 sky130_fd_sc_hd__nor2_1 _6141_ (.A(_2569_),
    .B(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__o21ai_1 _6142_ (.A1(_2483_),
    .A2(_2486_),
    .B1(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__or3_1 _6143_ (.A(_2483_),
    .B(_2486_),
    .C(_2571_),
    .X(_2573_));
 sky130_fd_sc_hd__or4bb_1 _6144_ (.A(_2525_),
    .B(_2526_),
    .C_N(_2572_),
    .D_N(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__a2bb2o_1 _6145_ (.A1_N(_2525_),
    .A2_N(_2526_),
    .B1(_2572_),
    .B2(_2573_),
    .X(_2575_));
 sky130_fd_sc_hd__and3_1 _6146_ (.A(_2507_),
    .B(_2574_),
    .C(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__a21o_1 _6147_ (.A1(_2574_),
    .A2(_2575_),
    .B1(_2507_),
    .X(_2577_));
 sky130_fd_sc_hd__nand2b_1 _6148_ (.A_N(_2576_),
    .B(_2577_),
    .Y(_2578_));
 sky130_fd_sc_hd__nor3b_1 _6149_ (.A(_2506_),
    .B(_2576_),
    .C_N(_2577_),
    .Y(_2579_));
 sky130_fd_sc_hd__and2_1 _6150_ (.A(_2506_),
    .B(_2578_),
    .X(_2580_));
 sky130_fd_sc_hd__or2_2 _6151_ (.A(_2579_),
    .B(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__and2b_1 _6152_ (.A_N(_2581_),
    .B(_2505_),
    .X(_2582_));
 sky130_fd_sc_hd__xnor2_1 _6153_ (.A(_2505_),
    .B(_2581_),
    .Y(_2583_));
 sky130_fd_sc_hd__xor2_1 _6154_ (.A(_2498_),
    .B(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__xnor2_1 _6155_ (.A(_2504_),
    .B(_2584_),
    .Y(_2585_));
 sky130_fd_sc_hd__nor2_1 _6156_ (.A(net194),
    .B(_2585_),
    .Y(_0021_));
 sky130_fd_sc_hd__o21a_1 _6157_ (.A1(_2498_),
    .A2(_2500_),
    .B1(_2583_),
    .X(_2586_));
 sky130_fd_sc_hd__a31o_1 _6158_ (.A1(_2421_),
    .A2(_2502_),
    .A3(_2584_),
    .B1(_2586_),
    .X(_2587_));
 sky130_fd_sc_hd__a21oi_1 _6159_ (.A1(_2522_),
    .A2(_2523_),
    .B1(_2525_),
    .Y(_2588_));
 sky130_fd_sc_hd__a21o_1 _6160_ (.A1(_2509_),
    .A2(_2518_),
    .B1(_2520_),
    .X(_2589_));
 sky130_fd_sc_hd__nand2_2 _6161_ (.A(_1360_),
    .B(_1536_),
    .Y(_2590_));
 sky130_fd_sc_hd__o21a_1 _6162_ (.A1(_1722_),
    .A2(_1821_),
    .B1(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__a21bo_1 _6163_ (.A1(_1725_),
    .A2(_2512_),
    .B1_N(_2511_),
    .X(_2592_));
 sky130_fd_sc_hd__and2b_1 _6164_ (.A_N(_2095_),
    .B(_1827_),
    .X(_2593_));
 sky130_fd_sc_hd__nand2b_1 _6165_ (.A_N(_2095_),
    .B(_1827_),
    .Y(_2594_));
 sky130_fd_sc_hd__and2b_1 _6166_ (.A_N(_1827_),
    .B(_2095_),
    .X(_2595_));
 sky130_fd_sc_hd__nor2_1 _6167_ (.A(_2593_),
    .B(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__xnor2_1 _6168_ (.A(_1822_),
    .B(_2596_),
    .Y(_2597_));
 sky130_fd_sc_hd__o21a_1 _6169_ (.A1(_2527_),
    .A2(_2530_),
    .B1(_2597_),
    .X(_2598_));
 sky130_fd_sc_hd__nor3_1 _6170_ (.A(_2527_),
    .B(_2530_),
    .C(_2597_),
    .Y(_2599_));
 sky130_fd_sc_hd__nor2_1 _6171_ (.A(_2598_),
    .B(_2599_),
    .Y(_2600_));
 sky130_fd_sc_hd__xor2_1 _6172_ (.A(_2592_),
    .B(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__o21a_1 _6173_ (.A1(_2514_),
    .A2(_2517_),
    .B1(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__nor3_1 _6174_ (.A(_2514_),
    .B(_2517_),
    .C(_2601_),
    .Y(_2603_));
 sky130_fd_sc_hd__nor2_1 _6175_ (.A(_2602_),
    .B(_2603_),
    .Y(_2604_));
 sky130_fd_sc_hd__and2_1 _6176_ (.A(_2591_),
    .B(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__nor2_1 _6177_ (.A(_2591_),
    .B(_2604_),
    .Y(_2606_));
 sky130_fd_sc_hd__or2_1 _6178_ (.A(_2605_),
    .B(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__a31oi_2 _6179_ (.A1(_2546_),
    .A2(_2547_),
    .A3(_2548_),
    .B1(_2552_),
    .Y(_2608_));
 sky130_fd_sc_hd__xnor2_1 _6180_ (.A(_2607_),
    .B(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__and2b_1 _6181_ (.A_N(_2609_),
    .B(_2589_),
    .X(_2610_));
 sky130_fd_sc_hd__xnor2_1 _6182_ (.A(_2589_),
    .B(_2609_),
    .Y(_2611_));
 sky130_fd_sc_hd__and2b_1 _6183_ (.A_N(_2362_),
    .B(_2367_),
    .X(_2612_));
 sky130_fd_sc_hd__and2b_1 _6184_ (.A_N(_2367_),
    .B(_2362_),
    .X(_2613_));
 sky130_fd_sc_hd__or2_1 _6185_ (.A(_2612_),
    .B(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__inv_2 _6186_ (.A(_2614_),
    .Y(_2615_));
 sky130_fd_sc_hd__xor2_2 _6187_ (.A(_2100_),
    .B(_2614_),
    .X(_2616_));
 sky130_fd_sc_hd__nand2_1 _6188_ (.A(_2540_),
    .B(_2542_),
    .Y(_2617_));
 sky130_fd_sc_hd__o21ai_1 _6189_ (.A1(net105),
    .A2(net108),
    .B1(net148),
    .Y(_2618_));
 sky130_fd_sc_hd__a21o_1 _6190_ (.A1(net105),
    .A2(net108),
    .B1(_2618_),
    .X(_2619_));
 sky130_fd_sc_hd__xnor2_1 _6191_ (.A(_2451_),
    .B(_2619_),
    .Y(_2620_));
 sky130_fd_sc_hd__o21ai_1 _6192_ (.A1(_2471_),
    .A2(_2555_),
    .B1(_2620_),
    .Y(_2621_));
 sky130_fd_sc_hd__or3_1 _6193_ (.A(_2471_),
    .B(_2555_),
    .C(_2620_),
    .X(_2622_));
 sky130_fd_sc_hd__a31o_1 _6194_ (.A1(net111),
    .A2(\ann.weight[15] ),
    .A3(_2536_),
    .B1(_2535_),
    .X(_2623_));
 sky130_fd_sc_hd__and3_1 _6195_ (.A(_2621_),
    .B(_2622_),
    .C(_2623_),
    .X(_2624_));
 sky130_fd_sc_hd__a21oi_1 _6196_ (.A1(_2621_),
    .A2(_2622_),
    .B1(_2623_),
    .Y(_2625_));
 sky130_fd_sc_hd__or2_1 _6197_ (.A(_2624_),
    .B(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__xnor2_1 _6198_ (.A(_2617_),
    .B(_2626_),
    .Y(_2627_));
 sky130_fd_sc_hd__nor2_1 _6199_ (.A(_2616_),
    .B(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__and2_1 _6200_ (.A(_2616_),
    .B(_2627_),
    .X(_2629_));
 sky130_fd_sc_hd__or2_1 _6201_ (.A(_2628_),
    .B(_2629_),
    .X(_2630_));
 sky130_fd_sc_hd__a21oi_1 _6202_ (.A1(_2558_),
    .A2(_2560_),
    .B1(_2630_),
    .Y(_2631_));
 sky130_fd_sc_hd__and3_1 _6203_ (.A(_2558_),
    .B(_2560_),
    .C(_2630_),
    .X(_2632_));
 sky130_fd_sc_hd__a211o_1 _6204_ (.A1(_2544_),
    .A2(_2546_),
    .B1(_2631_),
    .C1(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__o211ai_1 _6205_ (.A1(_2631_),
    .A2(_2632_),
    .B1(_2544_),
    .C1(_2546_),
    .Y(_2634_));
 sky130_fd_sc_hd__o21ai_1 _6206_ (.A1(_2391_),
    .A2(_2556_),
    .B1(_2383_),
    .Y(_2635_));
 sky130_fd_sc_hd__xor2_1 _6207_ (.A(_2559_),
    .B(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__xnor2_1 _6208_ (.A(_2228_),
    .B(_2636_),
    .Y(_2637_));
 sky130_fd_sc_hd__o21ba_1 _6209_ (.A1(_2227_),
    .A2(_2563_),
    .B1_N(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__or3b_1 _6210_ (.A(_2227_),
    .B(_2563_),
    .C_N(_2637_),
    .X(_2639_));
 sky130_fd_sc_hd__and2b_1 _6211_ (.A_N(_2638_),
    .B(_2639_),
    .X(_2640_));
 sky130_fd_sc_hd__and3_1 _6212_ (.A(_2633_),
    .B(_2634_),
    .C(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__a21oi_1 _6213_ (.A1(_2633_),
    .A2(_2634_),
    .B1(_2640_),
    .Y(_2642_));
 sky130_fd_sc_hd__nor2_1 _6214_ (.A(_2641_),
    .B(_2642_),
    .Y(_2643_));
 sky130_fd_sc_hd__o21ai_1 _6215_ (.A1(_2566_),
    .A2(_2569_),
    .B1(_2643_),
    .Y(_2644_));
 sky130_fd_sc_hd__or3_1 _6216_ (.A(_2566_),
    .B(_2569_),
    .C(_2643_),
    .X(_2645_));
 sky130_fd_sc_hd__nand2_1 _6217_ (.A(_2644_),
    .B(_2645_),
    .Y(_2646_));
 sky130_fd_sc_hd__xor2_1 _6218_ (.A(_2611_),
    .B(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__a21oi_1 _6219_ (.A1(_2572_),
    .A2(_2574_),
    .B1(_2647_),
    .Y(_2648_));
 sky130_fd_sc_hd__and3_1 _6220_ (.A(_2572_),
    .B(_2574_),
    .C(_2647_),
    .X(_2649_));
 sky130_fd_sc_hd__or3_1 _6221_ (.A(_2588_),
    .B(_2648_),
    .C(_2649_),
    .X(_2650_));
 sky130_fd_sc_hd__o21ai_1 _6222_ (.A1(_2648_),
    .A2(_2649_),
    .B1(_2588_),
    .Y(_2651_));
 sky130_fd_sc_hd__o211a_1 _6223_ (.A1(_2576_),
    .A2(_2579_),
    .B1(_2650_),
    .C1(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__a211o_1 _6224_ (.A1(_2650_),
    .A2(_2651_),
    .B1(_2576_),
    .C1(_2579_),
    .X(_2653_));
 sky130_fd_sc_hd__and2b_2 _6225_ (.A_N(_2652_),
    .B(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__and2_1 _6226_ (.A(_2582_),
    .B(_2654_),
    .X(_2655_));
 sky130_fd_sc_hd__nor2_1 _6227_ (.A(_2582_),
    .B(_2654_),
    .Y(_2656_));
 sky130_fd_sc_hd__nor2_1 _6228_ (.A(_2655_),
    .B(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__a21oi_1 _6229_ (.A1(_2587_),
    .A2(_2657_),
    .B1(net195),
    .Y(_2658_));
 sky130_fd_sc_hd__o21a_1 _6230_ (.A1(_2587_),
    .A2(_2657_),
    .B1(_2658_),
    .X(_0023_));
 sky130_fd_sc_hd__a21o_1 _6231_ (.A1(_2587_),
    .A2(_2657_),
    .B1(_2655_),
    .X(_2659_));
 sky130_fd_sc_hd__a21bo_1 _6232_ (.A1(_2559_),
    .A2(_2635_),
    .B1_N(_2558_),
    .X(_2660_));
 sky130_fd_sc_hd__and2b_1 _6233_ (.A_N(_2648_),
    .B(_2650_),
    .X(_2661_));
 sky130_fd_sc_hd__xor2_1 _6234_ (.A(_2652_),
    .B(_2661_),
    .X(_2662_));
 sky130_fd_sc_hd__mux2_1 _6235_ (.A0(_2621_),
    .A1(_2622_),
    .S(_2623_),
    .X(_2663_));
 sky130_fd_sc_hd__or4bb_1 _6236_ (.A(_2535_),
    .B(_2619_),
    .C_N(_2536_),
    .D_N(net148),
    .X(_2664_));
 sky130_fd_sc_hd__xnor2_1 _6237_ (.A(_2663_),
    .B(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__xnor2_1 _6238_ (.A(_2662_),
    .B(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__xnor2_2 _6239_ (.A(_2660_),
    .B(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__o21ba_1 _6240_ (.A1(_2607_),
    .A2(_2608_),
    .B1_N(_2610_),
    .X(_2668_));
 sky130_fd_sc_hd__xnor2_1 _6241_ (.A(_2590_),
    .B(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__a21oi_1 _6242_ (.A1(_2592_),
    .A2(_2600_),
    .B1(_2598_),
    .Y(_2670_));
 sky130_fd_sc_hd__and2b_1 _6243_ (.A_N(_2631_),
    .B(_2633_),
    .X(_2671_));
 sky130_fd_sc_hd__xnor2_1 _6244_ (.A(_2670_),
    .B(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__xnor2_1 _6245_ (.A(_2669_),
    .B(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__o21ai_1 _6246_ (.A1(_1822_),
    .A2(_2595_),
    .B1(_2594_),
    .Y(_2674_));
 sky130_fd_sc_hd__nor2_1 _6247_ (.A(_2602_),
    .B(_2605_),
    .Y(_2675_));
 sky130_fd_sc_hd__a21oi_1 _6248_ (.A1(_2100_),
    .A2(_2615_),
    .B1(_2612_),
    .Y(_2676_));
 sky130_fd_sc_hd__xnor2_1 _6249_ (.A(_2675_),
    .B(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__xnor2_1 _6250_ (.A(_2674_),
    .B(_2677_),
    .Y(_2678_));
 sky130_fd_sc_hd__xnor2_2 _6251_ (.A(_1911_),
    .B(_2678_),
    .Y(_2679_));
 sky130_fd_sc_hd__xnor2_2 _6252_ (.A(_2673_),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__xnor2_4 _6253_ (.A(_2667_),
    .B(_2680_),
    .Y(_2681_));
 sky130_fd_sc_hd__a221o_1 _6254_ (.A1(_0559_),
    .A2(_1536_),
    .B1(_1538_),
    .B2(_1359_),
    .C1(_1362_),
    .X(_2682_));
 sky130_fd_sc_hd__a21o_1 _6255_ (.A1(_2617_),
    .A2(_2626_),
    .B1(_2628_),
    .X(_2683_));
 sky130_fd_sc_hd__nor2_1 _6256_ (.A(_2638_),
    .B(_2641_),
    .Y(_2684_));
 sky130_fd_sc_hd__xnor2_2 _6257_ (.A(_2683_),
    .B(_2684_),
    .Y(_2685_));
 sky130_fd_sc_hd__xnor2_1 _6258_ (.A(_2682_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__xnor2_1 _6259_ (.A(_2190_),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__a21bo_1 _6260_ (.A1(_2611_),
    .A2(_2645_),
    .B1_N(_2644_),
    .X(_2688_));
 sky130_fd_sc_hd__xor2_1 _6261_ (.A(_2455_),
    .B(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__mux2_1 _6262_ (.A0(_2226_),
    .A1(_2227_),
    .S(_2636_),
    .X(_2690_));
 sky130_fd_sc_hd__xnor2_1 _6263_ (.A(_2689_),
    .B(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__xnor2_1 _6264_ (.A(_2687_),
    .B(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__xor2_1 _6265_ (.A(_2181_),
    .B(_2185_),
    .X(_2693_));
 sky130_fd_sc_hd__xnor2_1 _6266_ (.A(_2450_),
    .B(_2693_),
    .Y(_2694_));
 sky130_fd_sc_hd__xnor2_2 _6267_ (.A(_2692_),
    .B(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__xnor2_4 _6268_ (.A(_2681_),
    .B(_2695_),
    .Y(_2696_));
 sky130_fd_sc_hd__xnor2_1 _6269_ (.A(_2659_),
    .B(_2696_),
    .Y(_2697_));
 sky130_fd_sc_hd__nor2_1 _6270_ (.A(net194),
    .B(_2697_),
    .Y(_0024_));
 sky130_fd_sc_hd__and3_1 _6271_ (.A(\ann.X[0] ),
    .B(\ann.multiply_FF[0] ),
    .C(net201),
    .X(_2698_));
 sky130_fd_sc_hd__a21oi_1 _6272_ (.A1(\ann.multiply_FF[0] ),
    .A2(net201),
    .B1(\ann.X[0] ),
    .Y(_2699_));
 sky130_fd_sc_hd__or2_1 _6273_ (.A(\ann.bias[0] ),
    .B(\ann.sum[0] ),
    .X(_2700_));
 sky130_fd_sc_hd__nand2_1 _6274_ (.A(\ann.bias[0] ),
    .B(\ann.sum[0] ),
    .Y(_2701_));
 sky130_fd_sc_hd__o21ai_1 _6275_ (.A1(_2698_),
    .A2(_2699_),
    .B1(net67),
    .Y(_2702_));
 sky130_fd_sc_hd__a21o_1 _6276_ (.A1(_2700_),
    .A2(_2701_),
    .B1(net68),
    .X(_2703_));
 sky130_fd_sc_hd__and3_1 _6277_ (.A(net201),
    .B(_2702_),
    .C(_2703_),
    .X(_0032_));
 sky130_fd_sc_hd__a21o_1 _6278_ (.A1(\ann.multiply_FF[1] ),
    .A2(net202),
    .B1(\ann.X[1] ),
    .X(_2704_));
 sky130_fd_sc_hd__nand3_1 _6279_ (.A(\ann.X[1] ),
    .B(\ann.multiply_FF[1] ),
    .C(net201),
    .Y(_2705_));
 sky130_fd_sc_hd__a21oi_1 _6280_ (.A1(_2704_),
    .A2(_2705_),
    .B1(_2698_),
    .Y(_2706_));
 sky130_fd_sc_hd__and3_1 _6281_ (.A(_2698_),
    .B(_2704_),
    .C(_2705_),
    .X(_2707_));
 sky130_fd_sc_hd__and2_1 _6282_ (.A(\ann.bias[1] ),
    .B(\ann.sum[1] ),
    .X(_2708_));
 sky130_fd_sc_hd__xor2_1 _6283_ (.A(\ann.bias[1] ),
    .B(\ann.sum[1] ),
    .X(_2709_));
 sky130_fd_sc_hd__o21ai_1 _6284_ (.A1(_2706_),
    .A2(_2707_),
    .B1(net67),
    .Y(_2710_));
 sky130_fd_sc_hd__xnor2_1 _6285_ (.A(_2701_),
    .B(_2709_),
    .Y(_2711_));
 sky130_fd_sc_hd__o211a_1 _6286_ (.A1(net68),
    .A2(_2711_),
    .B1(_2710_),
    .C1(net201),
    .X(_0043_));
 sky130_fd_sc_hd__a21bo_1 _6287_ (.A1(_2698_),
    .A2(_2704_),
    .B1_N(_2705_),
    .X(_2712_));
 sky130_fd_sc_hd__a21o_1 _6288_ (.A1(\ann.multiply_FF[2] ),
    .A2(net203),
    .B1(\ann.X[2] ),
    .X(_2713_));
 sky130_fd_sc_hd__nand3_1 _6289_ (.A(\ann.X[2] ),
    .B(\ann.multiply_FF[2] ),
    .C(net203),
    .Y(_2714_));
 sky130_fd_sc_hd__and3_1 _6290_ (.A(_2712_),
    .B(_2713_),
    .C(_2714_),
    .X(_2715_));
 sky130_fd_sc_hd__a21oi_1 _6291_ (.A1(_2713_),
    .A2(_2714_),
    .B1(_2712_),
    .Y(_2716_));
 sky130_fd_sc_hd__o21ai_1 _6292_ (.A1(_2715_),
    .A2(_2716_),
    .B1(net68),
    .Y(_2717_));
 sky130_fd_sc_hd__a31oi_2 _6293_ (.A1(\ann.bias[0] ),
    .A2(\ann.sum[0] ),
    .A3(_2709_),
    .B1(_2708_),
    .Y(_2718_));
 sky130_fd_sc_hd__nor2_1 _6294_ (.A(\ann.bias[2] ),
    .B(\ann.sum[2] ),
    .Y(_2719_));
 sky130_fd_sc_hd__or2_1 _6295_ (.A(\ann.bias[2] ),
    .B(\ann.sum[2] ),
    .X(_2720_));
 sky130_fd_sc_hd__nand2_1 _6296_ (.A(\ann.bias[2] ),
    .B(\ann.sum[2] ),
    .Y(_2721_));
 sky130_fd_sc_hd__a21oi_1 _6297_ (.A1(_2720_),
    .A2(_2721_),
    .B1(_2718_),
    .Y(_2722_));
 sky130_fd_sc_hd__a31o_1 _6298_ (.A1(_2718_),
    .A2(_2720_),
    .A3(_2721_),
    .B1(net66),
    .X(_2723_));
 sky130_fd_sc_hd__o211a_1 _6299_ (.A1(_2722_),
    .A2(_2723_),
    .B1(net204),
    .C1(_2717_),
    .X(_0054_));
 sky130_fd_sc_hd__a21bo_1 _6300_ (.A1(_2712_),
    .A2(_2713_),
    .B1_N(_2714_),
    .X(_2724_));
 sky130_fd_sc_hd__a21o_1 _6301_ (.A1(\ann.multiply_FF[3] ),
    .A2(net203),
    .B1(\ann.X[3] ),
    .X(_2725_));
 sky130_fd_sc_hd__nand3_1 _6302_ (.A(\ann.X[3] ),
    .B(\ann.multiply_FF[3] ),
    .C(net203),
    .Y(_2726_));
 sky130_fd_sc_hd__nand2_1 _6303_ (.A(_2725_),
    .B(_2726_),
    .Y(_2727_));
 sky130_fd_sc_hd__xnor2_1 _6304_ (.A(_2724_),
    .B(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__o21a_1 _6305_ (.A1(_2718_),
    .A2(_2719_),
    .B1(_2721_),
    .X(_2729_));
 sky130_fd_sc_hd__nor2_1 _6306_ (.A(\ann.bias[3] ),
    .B(\ann.sum[3] ),
    .Y(_2730_));
 sky130_fd_sc_hd__nand2_1 _6307_ (.A(\ann.bias[3] ),
    .B(\ann.sum[3] ),
    .Y(_2731_));
 sky130_fd_sc_hd__and2b_1 _6308_ (.A_N(_2730_),
    .B(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__o21a_1 _6309_ (.A1(_2729_),
    .A2(_2732_),
    .B1(net62),
    .X(_2733_));
 sky130_fd_sc_hd__a21bo_1 _6310_ (.A1(_2729_),
    .A2(_2732_),
    .B1_N(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__o211a_1 _6311_ (.A1(net63),
    .A2(_2728_),
    .B1(_2734_),
    .C1(net203),
    .X(_0057_));
 sky130_fd_sc_hd__a21boi_1 _6312_ (.A1(_2724_),
    .A2(_2725_),
    .B1_N(_2726_),
    .Y(_2735_));
 sky130_fd_sc_hd__a21oi_1 _6313_ (.A1(\ann.multiply_FF[4] ),
    .A2(net203),
    .B1(\ann.X[4] ),
    .Y(_2736_));
 sky130_fd_sc_hd__and3_1 _6314_ (.A(\ann.X[4] ),
    .B(\ann.multiply_FF[4] ),
    .C(net203),
    .X(_2737_));
 sky130_fd_sc_hd__or2_1 _6315_ (.A(_2736_),
    .B(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__o21a_1 _6316_ (.A1(_2729_),
    .A2(_2730_),
    .B1(_2731_),
    .X(_2739_));
 sky130_fd_sc_hd__or2_1 _6317_ (.A(\ann.bias[4] ),
    .B(\ann.sum[4] ),
    .X(_2740_));
 sky130_fd_sc_hd__nand2_1 _6318_ (.A(\ann.bias[4] ),
    .B(\ann.sum[4] ),
    .Y(_2741_));
 sky130_fd_sc_hd__and2_1 _6319_ (.A(_2740_),
    .B(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__inv_2 _6320_ (.A(_2742_),
    .Y(_2743_));
 sky130_fd_sc_hd__xor2_1 _6321_ (.A(_2735_),
    .B(_2738_),
    .X(_2744_));
 sky130_fd_sc_hd__xnor2_1 _6322_ (.A(_2739_),
    .B(_2743_),
    .Y(_2745_));
 sky130_fd_sc_hd__nand2_1 _6323_ (.A(net62),
    .B(_2745_),
    .Y(_2746_));
 sky130_fd_sc_hd__o211a_1 _6324_ (.A1(net62),
    .A2(_2744_),
    .B1(_2746_),
    .C1(net203),
    .X(_0058_));
 sky130_fd_sc_hd__a21oi_2 _6325_ (.A1(\ann.multiply_FF[5] ),
    .A2(net203),
    .B1(\ann.X[5] ),
    .Y(_2747_));
 sky130_fd_sc_hd__nand3_2 _6326_ (.A(\ann.X[5] ),
    .B(\ann.multiply_FF[5] ),
    .C(net203),
    .Y(_2748_));
 sky130_fd_sc_hd__and2b_1 _6327_ (.A_N(_2747_),
    .B(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__o21ba_1 _6328_ (.A1(_2735_),
    .A2(_2738_),
    .B1_N(_2737_),
    .X(_2750_));
 sky130_fd_sc_hd__and2_1 _6329_ (.A(_2749_),
    .B(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__o21ai_1 _6330_ (.A1(_2749_),
    .A2(_2750_),
    .B1(net66),
    .Y(_2752_));
 sky130_fd_sc_hd__nor2_1 _6331_ (.A(\ann.bias[5] ),
    .B(\ann.sum[5] ),
    .Y(_2753_));
 sky130_fd_sc_hd__and2_1 _6332_ (.A(\ann.bias[5] ),
    .B(\ann.sum[5] ),
    .X(_2754_));
 sky130_fd_sc_hd__nor2_1 _6333_ (.A(_2753_),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__inv_2 _6334_ (.A(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__o21a_1 _6335_ (.A1(_2739_),
    .A2(_2743_),
    .B1(_2741_),
    .X(_2757_));
 sky130_fd_sc_hd__xnor2_1 _6336_ (.A(_2755_),
    .B(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__o221a_1 _6337_ (.A1(_2751_),
    .A2(_2752_),
    .B1(_2758_),
    .B2(net66),
    .C1(net203),
    .X(_0059_));
 sky130_fd_sc_hd__a21oi_2 _6338_ (.A1(\ann.multiply_FF[6] ),
    .A2(net203),
    .B1(\ann.X[6] ),
    .Y(_2759_));
 sky130_fd_sc_hd__and3_2 _6339_ (.A(\ann.X[6] ),
    .B(\ann.multiply_FF[6] ),
    .C(net203),
    .X(_2760_));
 sky130_fd_sc_hd__a21o_1 _6340_ (.A1(_2748_),
    .A2(_2750_),
    .B1(_2747_),
    .X(_2761_));
 sky130_fd_sc_hd__o21a_1 _6341_ (.A1(_2759_),
    .A2(_2760_),
    .B1(_2761_),
    .X(_2762_));
 sky130_fd_sc_hd__a2111oi_4 _6342_ (.A1(_2748_),
    .A2(_2750_),
    .B1(_2759_),
    .C1(_2760_),
    .D1(_2747_),
    .Y(_2763_));
 sky130_fd_sc_hd__or3_1 _6343_ (.A(net62),
    .B(_2762_),
    .C(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__or2_1 _6344_ (.A(\ann.bias[6] ),
    .B(\ann.sum[6] ),
    .X(_2765_));
 sky130_fd_sc_hd__nand2_1 _6345_ (.A(\ann.bias[6] ),
    .B(\ann.sum[6] ),
    .Y(_2766_));
 sky130_fd_sc_hd__nand2_1 _6346_ (.A(_2765_),
    .B(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__o211a_1 _6347_ (.A1(\ann.bias[5] ),
    .A2(\ann.sum[5] ),
    .B1(\ann.sum[4] ),
    .C1(\ann.bias[4] ),
    .X(_2768_));
 sky130_fd_sc_hd__nor2_1 _6348_ (.A(_2754_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__o31a_1 _6349_ (.A1(_2739_),
    .A2(_2743_),
    .A3(_2756_),
    .B1(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__and2_1 _6350_ (.A(_2767_),
    .B(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__or2_1 _6351_ (.A(_2767_),
    .B(_2770_),
    .X(_2772_));
 sky130_fd_sc_hd__or3b_1 _6352_ (.A(net67),
    .B(_2771_),
    .C_N(_2772_),
    .X(_2773_));
 sky130_fd_sc_hd__a21oi_1 _6353_ (.A1(_2764_),
    .A2(_2773_),
    .B1(net194),
    .Y(_0060_));
 sky130_fd_sc_hd__a21o_1 _6354_ (.A1(\ann.multiply_FF[7] ),
    .A2(net204),
    .B1(\ann.X[7] ),
    .X(_2774_));
 sky130_fd_sc_hd__nand3_1 _6355_ (.A(\ann.X[7] ),
    .B(\ann.multiply_FF[7] ),
    .C(net204),
    .Y(_2775_));
 sky130_fd_sc_hd__nand2_1 _6356_ (.A(_2774_),
    .B(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__o21ai_1 _6357_ (.A1(_2760_),
    .A2(_2763_),
    .B1(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__o31a_1 _6358_ (.A1(_2760_),
    .A2(_2763_),
    .A3(_2776_),
    .B1(net67),
    .X(_2778_));
 sky130_fd_sc_hd__nor2_1 _6359_ (.A(\ann.bias[7] ),
    .B(\ann.sum[7] ),
    .Y(_2779_));
 sky130_fd_sc_hd__nand2_1 _6360_ (.A(\ann.bias[7] ),
    .B(\ann.sum[7] ),
    .Y(_2780_));
 sky130_fd_sc_hd__and2b_1 _6361_ (.A_N(_2779_),
    .B(_2780_),
    .X(_2781_));
 sky130_fd_sc_hd__a21oi_1 _6362_ (.A1(_2766_),
    .A2(_2772_),
    .B1(_2781_),
    .Y(_2782_));
 sky130_fd_sc_hd__a31o_1 _6363_ (.A1(_2766_),
    .A2(_2772_),
    .A3(_2781_),
    .B1(net67),
    .X(_2783_));
 sky130_fd_sc_hd__o21ai_1 _6364_ (.A1(_2782_),
    .A2(_2783_),
    .B1(net204),
    .Y(_2784_));
 sky130_fd_sc_hd__a21oi_1 _6365_ (.A1(_2777_),
    .A2(_2778_),
    .B1(_2784_),
    .Y(_0061_));
 sky130_fd_sc_hd__a21oi_1 _6366_ (.A1(\ann.multiply_FF[8] ),
    .A2(net206),
    .B1(\ann.X[8] ),
    .Y(_2785_));
 sky130_fd_sc_hd__and3_1 _6367_ (.A(\ann.X[8] ),
    .B(\ann.multiply_FF[8] ),
    .C(net205),
    .X(_2786_));
 sky130_fd_sc_hd__nor2_1 _6368_ (.A(_2785_),
    .B(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__nand2b_1 _6369_ (.A_N(_2760_),
    .B(_2775_),
    .Y(_2788_));
 sky130_fd_sc_hd__o21a_1 _6370_ (.A1(_2763_),
    .A2(_2788_),
    .B1(_2774_),
    .X(_2789_));
 sky130_fd_sc_hd__nor2_1 _6371_ (.A(_2787_),
    .B(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__o211a_1 _6372_ (.A1(_2763_),
    .A2(_2788_),
    .B1(_2787_),
    .C1(_2774_),
    .X(_2791_));
 sky130_fd_sc_hd__or3_1 _6373_ (.A(net63),
    .B(_2790_),
    .C(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__or2_1 _6374_ (.A(\ann.bias[8] ),
    .B(\ann.sum[8] ),
    .X(_2793_));
 sky130_fd_sc_hd__nand2_2 _6375_ (.A(\ann.bias[8] ),
    .B(\ann.sum[8] ),
    .Y(_2794_));
 sky130_fd_sc_hd__nand2_1 _6376_ (.A(_2793_),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__o211a_1 _6377_ (.A1(_2767_),
    .A2(_2770_),
    .B1(_2780_),
    .C1(_2766_),
    .X(_2796_));
 sky130_fd_sc_hd__or2_1 _6378_ (.A(_2779_),
    .B(_2796_),
    .X(_2797_));
 sky130_fd_sc_hd__and2_1 _6379_ (.A(_2795_),
    .B(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__or2_1 _6380_ (.A(_2795_),
    .B(_2797_),
    .X(_2799_));
 sky130_fd_sc_hd__or3b_1 _6381_ (.A(net67),
    .B(_2798_),
    .C_N(_2799_),
    .X(_2800_));
 sky130_fd_sc_hd__a21oi_1 _6382_ (.A1(_2792_),
    .A2(_2800_),
    .B1(net195),
    .Y(_0062_));
 sky130_fd_sc_hd__a21oi_2 _6383_ (.A1(\ann.multiply_FF[9] ),
    .A2(net206),
    .B1(\ann.X[9] ),
    .Y(_2801_));
 sky130_fd_sc_hd__inv_2 _6384_ (.A(_2801_),
    .Y(_2802_));
 sky130_fd_sc_hd__and3_1 _6385_ (.A(\ann.X[9] ),
    .B(\ann.multiply_FF[9] ),
    .C(net205),
    .X(_2803_));
 sky130_fd_sc_hd__o22a_1 _6386_ (.A1(_2786_),
    .A2(_2791_),
    .B1(_2801_),
    .B2(_2803_),
    .X(_2804_));
 sky130_fd_sc_hd__nor4_1 _6387_ (.A(_2786_),
    .B(_2791_),
    .C(_2801_),
    .D(_2803_),
    .Y(_2805_));
 sky130_fd_sc_hd__or2_2 _6388_ (.A(\ann.bias[9] ),
    .B(\ann.sum[9] ),
    .X(_2806_));
 sky130_fd_sc_hd__nand2_1 _6389_ (.A(\ann.bias[9] ),
    .B(\ann.sum[9] ),
    .Y(_2807_));
 sky130_fd_sc_hd__and4_1 _6390_ (.A(_2794_),
    .B(_2799_),
    .C(_2806_),
    .D(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__a22o_1 _6391_ (.A1(_2794_),
    .A2(_2799_),
    .B1(_2806_),
    .B2(_2807_),
    .X(_2809_));
 sky130_fd_sc_hd__or3b_1 _6392_ (.A(net67),
    .B(_2808_),
    .C_N(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__o311a_1 _6393_ (.A1(net63),
    .A2(_2804_),
    .A3(_2805_),
    .B1(_2810_),
    .C1(net205),
    .X(_0063_));
 sky130_fd_sc_hd__a21oi_1 _6394_ (.A1(\ann.multiply_FF[10] ),
    .A2(net205),
    .B1(\ann.X[10] ),
    .Y(_2811_));
 sky130_fd_sc_hd__and3_1 _6395_ (.A(\ann.X[10] ),
    .B(\ann.multiply_FF[10] ),
    .C(net205),
    .X(_2812_));
 sky130_fd_sc_hd__nor2_1 _6396_ (.A(_2811_),
    .B(_2812_),
    .Y(_2813_));
 sky130_fd_sc_hd__or2_1 _6397_ (.A(_2786_),
    .B(_2803_),
    .X(_2814_));
 sky130_fd_sc_hd__o21a_1 _6398_ (.A1(_2791_),
    .A2(_2814_),
    .B1(_2802_),
    .X(_2815_));
 sky130_fd_sc_hd__nor2_1 _6399_ (.A(_2813_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__o211a_1 _6400_ (.A1(_2791_),
    .A2(_2814_),
    .B1(_2813_),
    .C1(_2802_),
    .X(_2817_));
 sky130_fd_sc_hd__or3_1 _6401_ (.A(net63),
    .B(_2816_),
    .C(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__and2_1 _6402_ (.A(\ann.bias[10] ),
    .B(\ann.sum[10] ),
    .X(_2819_));
 sky130_fd_sc_hd__nand2_1 _6403_ (.A(\ann.bias[10] ),
    .B(\ann.sum[10] ),
    .Y(_2820_));
 sky130_fd_sc_hd__or2_1 _6404_ (.A(\ann.bias[10] ),
    .B(\ann.sum[10] ),
    .X(_2821_));
 sky130_fd_sc_hd__o311ai_4 _6405_ (.A1(_2779_),
    .A2(_2795_),
    .A3(_2796_),
    .B1(_2807_),
    .C1(_2794_),
    .Y(_2822_));
 sky130_fd_sc_hd__a22o_1 _6406_ (.A1(_2820_),
    .A2(_2821_),
    .B1(_2822_),
    .B2(_2806_),
    .X(_2823_));
 sky130_fd_sc_hd__nand4_1 _6407_ (.A(_2806_),
    .B(_2820_),
    .C(_2821_),
    .D(_2822_),
    .Y(_2824_));
 sky130_fd_sc_hd__nand3_1 _6408_ (.A(net63),
    .B(_2823_),
    .C(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__a21oi_1 _6409_ (.A1(_2818_),
    .A2(_2825_),
    .B1(net194),
    .Y(_0033_));
 sky130_fd_sc_hd__a21o_1 _6410_ (.A1(\ann.multiply_FF[11] ),
    .A2(net205),
    .B1(\ann.X[11] ),
    .X(_2826_));
 sky130_fd_sc_hd__nand3_2 _6411_ (.A(\ann.X[11] ),
    .B(\ann.multiply_FF[11] ),
    .C(net205),
    .Y(_2827_));
 sky130_fd_sc_hd__a211o_1 _6412_ (.A1(_2826_),
    .A2(_2827_),
    .B1(_2812_),
    .C1(_2817_),
    .X(_2828_));
 sky130_fd_sc_hd__o211ai_2 _6413_ (.A1(_2812_),
    .A2(_2817_),
    .B1(_2826_),
    .C1(_2827_),
    .Y(_2829_));
 sky130_fd_sc_hd__a31o_1 _6414_ (.A1(_2806_),
    .A2(_2821_),
    .A3(_2822_),
    .B1(_2819_),
    .X(_2830_));
 sky130_fd_sc_hd__nand2_1 _6415_ (.A(\ann.bias[11] ),
    .B(\ann.sum[11] ),
    .Y(_2831_));
 sky130_fd_sc_hd__or2_1 _6416_ (.A(\ann.bias[11] ),
    .B(\ann.sum[11] ),
    .X(_2832_));
 sky130_fd_sc_hd__nand2_1 _6417_ (.A(_2831_),
    .B(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__a21o_1 _6418_ (.A1(_2828_),
    .A2(_2829_),
    .B1(net63),
    .X(_2834_));
 sky130_fd_sc_hd__xnor2_1 _6419_ (.A(_2830_),
    .B(_2833_),
    .Y(_2835_));
 sky130_fd_sc_hd__o211a_1 _6420_ (.A1(net68),
    .A2(_2835_),
    .B1(_2834_),
    .C1(net206),
    .X(_0034_));
 sky130_fd_sc_hd__a21oi_1 _6421_ (.A1(\ann.multiply_FF[12] ),
    .A2(net205),
    .B1(\ann.X[12] ),
    .Y(_2836_));
 sky130_fd_sc_hd__and3_1 _6422_ (.A(\ann.X[12] ),
    .B(\ann.multiply_FF[12] ),
    .C(net205),
    .X(_2837_));
 sky130_fd_sc_hd__nand3_1 _6423_ (.A(\ann.X[12] ),
    .B(\ann.multiply_FF[12] ),
    .C(net205),
    .Y(_2838_));
 sky130_fd_sc_hd__o211ai_1 _6424_ (.A1(_2836_),
    .A2(_2837_),
    .B1(_2827_),
    .C1(_2829_),
    .Y(_2839_));
 sky130_fd_sc_hd__a211o_1 _6425_ (.A1(_2827_),
    .A2(_2829_),
    .B1(_2836_),
    .C1(_2837_),
    .X(_2840_));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(\ann.bias[12] ),
    .B(\ann.sum[12] ),
    .Y(_2841_));
 sky130_fd_sc_hd__or2_1 _6427_ (.A(\ann.bias[12] ),
    .B(\ann.sum[12] ),
    .X(_2842_));
 sky130_fd_sc_hd__a21bo_1 _6428_ (.A1(_2830_),
    .A2(_2832_),
    .B1_N(_2831_),
    .X(_2843_));
 sky130_fd_sc_hd__a21o_1 _6429_ (.A1(_2841_),
    .A2(_2842_),
    .B1(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__a31oi_1 _6430_ (.A1(_2841_),
    .A2(_2842_),
    .A3(_2843_),
    .B1(net68),
    .Y(_2845_));
 sky130_fd_sc_hd__a32o_1 _6431_ (.A1(net68),
    .A2(_2839_),
    .A3(_2840_),
    .B1(_2844_),
    .B2(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__and2_1 _6432_ (.A(net206),
    .B(_2846_),
    .X(_0035_));
 sky130_fd_sc_hd__a21oi_1 _6433_ (.A1(\ann.multiply_FF[13] ),
    .A2(net206),
    .B1(\ann.X[13] ),
    .Y(_2847_));
 sky130_fd_sc_hd__and3_1 _6434_ (.A(\ann.X[13] ),
    .B(\ann.multiply_FF[13] ),
    .C(net206),
    .X(_2848_));
 sky130_fd_sc_hd__nand3_1 _6435_ (.A(\ann.X[13] ),
    .B(\ann.multiply_FF[13] ),
    .C(net207),
    .Y(_2849_));
 sky130_fd_sc_hd__o211ai_1 _6436_ (.A1(_2847_),
    .A2(_2848_),
    .B1(_2838_),
    .C1(_2840_),
    .Y(_2850_));
 sky130_fd_sc_hd__a211o_1 _6437_ (.A1(_2838_),
    .A2(_2840_),
    .B1(_2847_),
    .C1(_2848_),
    .X(_2851_));
 sky130_fd_sc_hd__a21bo_1 _6438_ (.A1(_2842_),
    .A2(_2843_),
    .B1_N(_2841_),
    .X(_2852_));
 sky130_fd_sc_hd__nand2_1 _6439_ (.A(\ann.bias[13] ),
    .B(\ann.sum[13] ),
    .Y(_2853_));
 sky130_fd_sc_hd__or2_1 _6440_ (.A(\ann.bias[13] ),
    .B(\ann.sum[13] ),
    .X(_2854_));
 sky130_fd_sc_hd__nand2_1 _6441_ (.A(_2853_),
    .B(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__a21o_1 _6442_ (.A1(_2850_),
    .A2(_2851_),
    .B1(net63),
    .X(_2856_));
 sky130_fd_sc_hd__xnor2_1 _6443_ (.A(_2852_),
    .B(_2855_),
    .Y(_2857_));
 sky130_fd_sc_hd__o211a_1 _6444_ (.A1(net67),
    .A2(_2857_),
    .B1(_2856_),
    .C1(net206),
    .X(_0036_));
 sky130_fd_sc_hd__a21oi_1 _6445_ (.A1(\ann.multiply_FF[14] ),
    .A2(net207),
    .B1(\ann.X[14] ),
    .Y(_2858_));
 sky130_fd_sc_hd__and3_1 _6446_ (.A(\ann.X[14] ),
    .B(\ann.multiply_FF[14] ),
    .C(net207),
    .X(_2859_));
 sky130_fd_sc_hd__nand3_1 _6447_ (.A(\ann.X[14] ),
    .B(\ann.multiply_FF[14] ),
    .C(net202),
    .Y(_2860_));
 sky130_fd_sc_hd__o211a_1 _6448_ (.A1(_2858_),
    .A2(_2859_),
    .B1(_2849_),
    .C1(_2851_),
    .X(_2861_));
 sky130_fd_sc_hd__a211o_1 _6449_ (.A1(_2849_),
    .A2(_2851_),
    .B1(_2858_),
    .C1(_2859_),
    .X(_2862_));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(net68),
    .B(_2862_),
    .Y(_2863_));
 sky130_fd_sc_hd__nand2_1 _6451_ (.A(\ann.bias[14] ),
    .B(\ann.sum[14] ),
    .Y(_2864_));
 sky130_fd_sc_hd__or2_1 _6452_ (.A(\ann.bias[14] ),
    .B(\ann.sum[14] ),
    .X(_2865_));
 sky130_fd_sc_hd__nand2_1 _6453_ (.A(_2864_),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__a21boi_1 _6454_ (.A1(_2852_),
    .A2(_2854_),
    .B1_N(_2853_),
    .Y(_2867_));
 sky130_fd_sc_hd__and2_1 _6455_ (.A(_2866_),
    .B(_2867_),
    .X(_2868_));
 sky130_fd_sc_hd__nor2_1 _6456_ (.A(_2866_),
    .B(_2867_),
    .Y(_2869_));
 sky130_fd_sc_hd__o32a_1 _6457_ (.A1(net68),
    .A2(_2868_),
    .A3(_2869_),
    .B1(_2861_),
    .B2(_2863_),
    .X(_2870_));
 sky130_fd_sc_hd__nor2_1 _6458_ (.A(net194),
    .B(_2870_),
    .Y(_0037_));
 sky130_fd_sc_hd__a21oi_1 _6459_ (.A1(\ann.multiply_FF[15] ),
    .A2(net202),
    .B1(\ann.X[15] ),
    .Y(_2871_));
 sky130_fd_sc_hd__and3_1 _6460_ (.A(\ann.X[15] ),
    .B(\ann.multiply_FF[15] ),
    .C(net202),
    .X(_2872_));
 sky130_fd_sc_hd__o211a_1 _6461_ (.A1(_2871_),
    .A2(_2872_),
    .B1(_2860_),
    .C1(_2862_),
    .X(_2873_));
 sky130_fd_sc_hd__a211oi_2 _6462_ (.A1(_2860_),
    .A2(_2862_),
    .B1(_2871_),
    .C1(_2872_),
    .Y(_2874_));
 sky130_fd_sc_hd__o21a_1 _6463_ (.A1(_2866_),
    .A2(_2867_),
    .B1(_2864_),
    .X(_2875_));
 sky130_fd_sc_hd__nand2_1 _6464_ (.A(\ann.bias[15] ),
    .B(\ann.sum[15] ),
    .Y(_2876_));
 sky130_fd_sc_hd__or2_1 _6465_ (.A(\ann.bias[15] ),
    .B(\ann.sum[15] ),
    .X(_2877_));
 sky130_fd_sc_hd__nand2_1 _6466_ (.A(_2876_),
    .B(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__nand2_1 _6467_ (.A(_2875_),
    .B(_2878_),
    .Y(_2879_));
 sky130_fd_sc_hd__or2_1 _6468_ (.A(_2875_),
    .B(_2878_),
    .X(_2880_));
 sky130_fd_sc_hd__o21ai_1 _6469_ (.A1(_2873_),
    .A2(_2874_),
    .B1(net67),
    .Y(_2881_));
 sky130_fd_sc_hd__a21o_1 _6470_ (.A1(_2879_),
    .A2(_2880_),
    .B1(net68),
    .X(_2882_));
 sky130_fd_sc_hd__and3_1 _6471_ (.A(net202),
    .B(_2881_),
    .C(_2882_),
    .X(_0038_));
 sky130_fd_sc_hd__a21oi_1 _6472_ (.A1(\ann.multiply_FF[16] ),
    .A2(net201),
    .B1(\ann.X[16] ),
    .Y(_2883_));
 sky130_fd_sc_hd__and3_1 _6473_ (.A(\ann.X[16] ),
    .B(\ann.multiply_FF[16] ),
    .C(net201),
    .X(_2884_));
 sky130_fd_sc_hd__nor2_1 _6474_ (.A(_2883_),
    .B(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__or3_1 _6475_ (.A(_2872_),
    .B(_2874_),
    .C(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__o21a_1 _6476_ (.A1(_2872_),
    .A2(_2874_),
    .B1(_2885_),
    .X(_2887_));
 sky130_fd_sc_hd__or3b_1 _6477_ (.A(_2887_),
    .B(net63),
    .C_N(_2886_),
    .X(_2888_));
 sky130_fd_sc_hd__o21ai_2 _6478_ (.A1(_2875_),
    .A2(_2878_),
    .B1(_2876_),
    .Y(_2889_));
 sky130_fd_sc_hd__xnor2_1 _6479_ (.A(\ann.bias[16] ),
    .B(\ann.sum[16] ),
    .Y(_2890_));
 sky130_fd_sc_hd__inv_2 _6480_ (.A(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__nor2_1 _6481_ (.A(_2889_),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__and2_1 _6482_ (.A(_2889_),
    .B(_2891_),
    .X(_2893_));
 sky130_fd_sc_hd__or3_1 _6483_ (.A(net68),
    .B(_2892_),
    .C(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__a21oi_1 _6484_ (.A1(_2888_),
    .A2(_2894_),
    .B1(net194),
    .Y(_0039_));
 sky130_fd_sc_hd__a21oi_2 _6485_ (.A1(\ann.multiply_FF[17] ),
    .A2(net201),
    .B1(\ann.X[17] ),
    .Y(_2895_));
 sky130_fd_sc_hd__inv_2 _6486_ (.A(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__and3_1 _6487_ (.A(\ann.X[17] ),
    .B(\ann.multiply_FF[17] ),
    .C(net201),
    .X(_2897_));
 sky130_fd_sc_hd__o22a_1 _6488_ (.A1(_2884_),
    .A2(_2887_),
    .B1(_2895_),
    .B2(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__nor4_1 _6489_ (.A(_2884_),
    .B(_2887_),
    .C(_2895_),
    .D(_2897_),
    .Y(_2899_));
 sky130_fd_sc_hd__nor2_1 _6490_ (.A(\ann.bias[17] ),
    .B(\ann.sum[17] ),
    .Y(_2900_));
 sky130_fd_sc_hd__or2_1 _6491_ (.A(\ann.bias[17] ),
    .B(\ann.sum[17] ),
    .X(_2901_));
 sky130_fd_sc_hd__and2_1 _6492_ (.A(\ann.bias[17] ),
    .B(\ann.sum[17] ),
    .X(_2902_));
 sky130_fd_sc_hd__nor2_1 _6493_ (.A(_2900_),
    .B(_2902_),
    .Y(_2903_));
 sky130_fd_sc_hd__a21oi_1 _6494_ (.A1(\ann.bias[16] ),
    .A2(\ann.sum[16] ),
    .B1(_2893_),
    .Y(_2904_));
 sky130_fd_sc_hd__xnor2_1 _6495_ (.A(_2903_),
    .B(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__or2_1 _6496_ (.A(net66),
    .B(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__o311a_1 _6497_ (.A1(net62),
    .A2(_2898_),
    .A3(_2899_),
    .B1(_2906_),
    .C1(net201),
    .X(_0040_));
 sky130_fd_sc_hd__a21oi_1 _6498_ (.A1(\ann.multiply_FF[18] ),
    .A2(net202),
    .B1(\ann.X[18] ),
    .Y(_2907_));
 sky130_fd_sc_hd__and3_1 _6499_ (.A(\ann.X[18] ),
    .B(\ann.multiply_FF[18] ),
    .C(net202),
    .X(_2908_));
 sky130_fd_sc_hd__nor2_1 _6500_ (.A(_2907_),
    .B(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__or2_1 _6501_ (.A(_2884_),
    .B(_2897_),
    .X(_2910_));
 sky130_fd_sc_hd__or2_1 _6502_ (.A(_2887_),
    .B(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__a21oi_1 _6503_ (.A1(_2896_),
    .A2(_2911_),
    .B1(_2909_),
    .Y(_2912_));
 sky130_fd_sc_hd__o211a_1 _6504_ (.A1(_2887_),
    .A2(_2910_),
    .B1(_2909_),
    .C1(_2896_),
    .X(_2913_));
 sky130_fd_sc_hd__nand2_1 _6505_ (.A(\ann.bias[18] ),
    .B(\ann.sum[18] ),
    .Y(_2914_));
 sky130_fd_sc_hd__or2_1 _6506_ (.A(\ann.bias[18] ),
    .B(\ann.sum[18] ),
    .X(_2915_));
 sky130_fd_sc_hd__nand2_1 _6507_ (.A(_2914_),
    .B(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__a31o_1 _6508_ (.A1(\ann.bias[16] ),
    .A2(\ann.sum[16] ),
    .A3(_2901_),
    .B1(_2902_),
    .X(_2917_));
 sky130_fd_sc_hd__a31o_1 _6509_ (.A1(_2889_),
    .A2(_2891_),
    .A3(_2903_),
    .B1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__o21ai_1 _6510_ (.A1(_2912_),
    .A2(_2913_),
    .B1(net67),
    .Y(_2919_));
 sky130_fd_sc_hd__xnor2_1 _6511_ (.A(_2916_),
    .B(_2918_),
    .Y(_2920_));
 sky130_fd_sc_hd__o211a_1 _6512_ (.A1(net66),
    .A2(_2920_),
    .B1(_2919_),
    .C1(net204),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _6513_ (.A1(\ann.multiply_FF[19] ),
    .A2(net199),
    .B1(\ann.X[19] ),
    .X(_2921_));
 sky130_fd_sc_hd__nand3_1 _6514_ (.A(\ann.X[19] ),
    .B(\ann.multiply_FF[19] ),
    .C(net199),
    .Y(_2922_));
 sky130_fd_sc_hd__and2_1 _6515_ (.A(_2921_),
    .B(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__or3_1 _6516_ (.A(_2908_),
    .B(_2913_),
    .C(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__o21ai_2 _6517_ (.A1(_2908_),
    .A2(_2913_),
    .B1(_2923_),
    .Y(_2925_));
 sky130_fd_sc_hd__a21bo_1 _6518_ (.A1(_2915_),
    .A2(_2918_),
    .B1_N(_2914_),
    .X(_2926_));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(\ann.bias[19] ),
    .B(\ann.sum[19] ),
    .Y(_2927_));
 sky130_fd_sc_hd__or2_1 _6520_ (.A(\ann.bias[19] ),
    .B(\ann.sum[19] ),
    .X(_2928_));
 sky130_fd_sc_hd__a21o_1 _6521_ (.A1(_2927_),
    .A2(_2928_),
    .B1(_2926_),
    .X(_2929_));
 sky130_fd_sc_hd__a31oi_1 _6522_ (.A1(_2926_),
    .A2(_2927_),
    .A3(_2928_),
    .B1(net66),
    .Y(_2930_));
 sky130_fd_sc_hd__a32o_1 _6523_ (.A1(net67),
    .A2(_2924_),
    .A3(_2925_),
    .B1(_2929_),
    .B2(_2930_),
    .X(_2931_));
 sky130_fd_sc_hd__and2_1 _6524_ (.A(net199),
    .B(_2931_),
    .X(_0042_));
 sky130_fd_sc_hd__a21oi_1 _6525_ (.A1(\ann.multiply_FF[20] ),
    .A2(net199),
    .B1(\ann.X[20] ),
    .Y(_2932_));
 sky130_fd_sc_hd__and3_1 _6526_ (.A(\ann.X[20] ),
    .B(\ann.multiply_FF[20] ),
    .C(net199),
    .X(_2933_));
 sky130_fd_sc_hd__o211a_1 _6527_ (.A1(_2932_),
    .A2(_2933_),
    .B1(_2922_),
    .C1(_2925_),
    .X(_2934_));
 sky130_fd_sc_hd__a211oi_2 _6528_ (.A1(_2922_),
    .A2(_2925_),
    .B1(_2932_),
    .C1(_2933_),
    .Y(_2935_));
 sky130_fd_sc_hd__nand2_1 _6529_ (.A(\ann.bias[20] ),
    .B(\ann.sum[20] ),
    .Y(_2936_));
 sky130_fd_sc_hd__or2_1 _6530_ (.A(\ann.bias[20] ),
    .B(\ann.sum[20] ),
    .X(_2937_));
 sky130_fd_sc_hd__nand2_1 _6531_ (.A(_2936_),
    .B(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__a21bo_1 _6532_ (.A1(_2926_),
    .A2(_2928_),
    .B1_N(_2927_),
    .X(_2939_));
 sky130_fd_sc_hd__o21ai_1 _6533_ (.A1(_2934_),
    .A2(_2935_),
    .B1(net67),
    .Y(_2940_));
 sky130_fd_sc_hd__xnor2_1 _6534_ (.A(_2938_),
    .B(_2939_),
    .Y(_2941_));
 sky130_fd_sc_hd__o211a_1 _6535_ (.A1(net66),
    .A2(_2941_),
    .B1(_2940_),
    .C1(net197),
    .X(_0044_));
 sky130_fd_sc_hd__a21o_1 _6536_ (.A1(\ann.multiply_FF[21] ),
    .A2(net200),
    .B1(\ann.X[21] ),
    .X(_2942_));
 sky130_fd_sc_hd__nand3_2 _6537_ (.A(\ann.X[21] ),
    .B(\ann.multiply_FF[21] ),
    .C(net200),
    .Y(_2943_));
 sky130_fd_sc_hd__and2_1 _6538_ (.A(_2942_),
    .B(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__or3_1 _6539_ (.A(_2933_),
    .B(_2935_),
    .C(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__o21ai_2 _6540_ (.A1(_2933_),
    .A2(_2935_),
    .B1(_2944_),
    .Y(_2946_));
 sky130_fd_sc_hd__a21bo_1 _6541_ (.A1(_2937_),
    .A2(_2939_),
    .B1_N(_2936_),
    .X(_2947_));
 sky130_fd_sc_hd__nand2_1 _6542_ (.A(\ann.bias[21] ),
    .B(\ann.sum[21] ),
    .Y(_2948_));
 sky130_fd_sc_hd__or2_1 _6543_ (.A(\ann.bias[21] ),
    .B(\ann.sum[21] ),
    .X(_2949_));
 sky130_fd_sc_hd__a21o_1 _6544_ (.A1(_2948_),
    .A2(_2949_),
    .B1(_2947_),
    .X(_2950_));
 sky130_fd_sc_hd__a31oi_1 _6545_ (.A1(_2947_),
    .A2(_2948_),
    .A3(_2949_),
    .B1(net66),
    .Y(_2951_));
 sky130_fd_sc_hd__a32o_1 _6546_ (.A1(net66),
    .A2(_2945_),
    .A3(_2946_),
    .B1(_2950_),
    .B2(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__and2_1 _6547_ (.A(net197),
    .B(_2952_),
    .X(_0045_));
 sky130_fd_sc_hd__a21oi_2 _6548_ (.A1(\ann.multiply_FF[22] ),
    .A2(net200),
    .B1(\ann.X[22] ),
    .Y(_2953_));
 sky130_fd_sc_hd__and3_4 _6549_ (.A(\ann.X[22] ),
    .B(\ann.multiply_FF[22] ),
    .C(net200),
    .X(_2954_));
 sky130_fd_sc_hd__o211a_1 _6550_ (.A1(_2953_),
    .A2(_2954_),
    .B1(_2943_),
    .C1(_2946_),
    .X(_2955_));
 sky130_fd_sc_hd__a211oi_4 _6551_ (.A1(_2943_),
    .A2(_2946_),
    .B1(_2953_),
    .C1(_2954_),
    .Y(_2956_));
 sky130_fd_sc_hd__nand2_1 _6552_ (.A(\ann.bias[22] ),
    .B(\ann.sum[22] ),
    .Y(_2957_));
 sky130_fd_sc_hd__or2_1 _6553_ (.A(\ann.bias[22] ),
    .B(\ann.sum[22] ),
    .X(_2958_));
 sky130_fd_sc_hd__nand2_1 _6554_ (.A(_2957_),
    .B(_2958_),
    .Y(_2959_));
 sky130_fd_sc_hd__a21bo_1 _6555_ (.A1(_2947_),
    .A2(_2949_),
    .B1_N(_2948_),
    .X(_2960_));
 sky130_fd_sc_hd__o21ai_1 _6556_ (.A1(_2955_),
    .A2(_2956_),
    .B1(net66),
    .Y(_2961_));
 sky130_fd_sc_hd__xnor2_1 _6557_ (.A(_2959_),
    .B(_2960_),
    .Y(_2962_));
 sky130_fd_sc_hd__o211a_1 _6558_ (.A1(net66),
    .A2(_2962_),
    .B1(_2961_),
    .C1(net197),
    .X(_0046_));
 sky130_fd_sc_hd__nor2_1 _6559_ (.A(_2954_),
    .B(_2956_),
    .Y(_2963_));
 sky130_fd_sc_hd__a21o_2 _6560_ (.A1(\ann.multiply_FF[23] ),
    .A2(net197),
    .B1(\ann.X[23] ),
    .X(_2964_));
 sky130_fd_sc_hd__and3_2 _6561_ (.A(\ann.X[23] ),
    .B(\ann.multiply_FF[23] ),
    .C(net197),
    .X(_2965_));
 sky130_fd_sc_hd__inv_2 _6562_ (.A(_2965_),
    .Y(_2966_));
 sky130_fd_sc_hd__a21oi_1 _6563_ (.A1(_2964_),
    .A2(_2966_),
    .B1(_2963_),
    .Y(_2967_));
 sky130_fd_sc_hd__a31o_1 _6564_ (.A1(_2963_),
    .A2(_2964_),
    .A3(_2966_),
    .B1(net62),
    .X(_2968_));
 sky130_fd_sc_hd__a21bo_1 _6565_ (.A1(_2958_),
    .A2(_2960_),
    .B1_N(_2957_),
    .X(_2969_));
 sky130_fd_sc_hd__nand2_1 _6566_ (.A(\ann.bias[23] ),
    .B(\ann.sum[23] ),
    .Y(_2970_));
 sky130_fd_sc_hd__or2_1 _6567_ (.A(\ann.bias[23] ),
    .B(\ann.sum[23] ),
    .X(_2971_));
 sky130_fd_sc_hd__nand2_1 _6568_ (.A(_2970_),
    .B(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__xor2_1 _6569_ (.A(_2969_),
    .B(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__nand2_1 _6570_ (.A(net62),
    .B(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__o211a_1 _6571_ (.A1(_2967_),
    .A2(_2968_),
    .B1(_2974_),
    .C1(net197),
    .X(_0047_));
 sky130_fd_sc_hd__o31a_1 _6572_ (.A1(_2954_),
    .A2(_2956_),
    .A3(_2965_),
    .B1(_2964_),
    .X(_2975_));
 sky130_fd_sc_hd__nand3_1 _6573_ (.A(\ann.X[24] ),
    .B(\ann.multiply_FF[24] ),
    .C(net196),
    .Y(_2976_));
 sky130_fd_sc_hd__inv_2 _6574_ (.A(_2976_),
    .Y(_2977_));
 sky130_fd_sc_hd__a21oi_1 _6575_ (.A1(\ann.multiply_FF[24] ),
    .A2(net196),
    .B1(\ann.X[24] ),
    .Y(_2978_));
 sky130_fd_sc_hd__nor2_1 _6576_ (.A(_2977_),
    .B(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__nor2_1 _6577_ (.A(_2975_),
    .B(_2979_),
    .Y(_2980_));
 sky130_fd_sc_hd__o311a_1 _6578_ (.A1(_2954_),
    .A2(_2956_),
    .A3(_2965_),
    .B1(_2979_),
    .C1(_2964_),
    .X(_2981_));
 sky130_fd_sc_hd__a21bo_1 _6579_ (.A1(_2969_),
    .A2(_2971_),
    .B1_N(_2970_),
    .X(_2982_));
 sky130_fd_sc_hd__and2_1 _6580_ (.A(\ann.bias[24] ),
    .B(\ann.sum[24] ),
    .X(_2983_));
 sky130_fd_sc_hd__nor2_1 _6581_ (.A(\ann.bias[24] ),
    .B(\ann.sum[24] ),
    .Y(_2984_));
 sky130_fd_sc_hd__nor2_1 _6582_ (.A(_2983_),
    .B(_2984_),
    .Y(_2985_));
 sky130_fd_sc_hd__o21ai_1 _6583_ (.A1(_2980_),
    .A2(_2981_),
    .B1(net66),
    .Y(_2986_));
 sky130_fd_sc_hd__xor2_1 _6584_ (.A(_2982_),
    .B(_2985_),
    .X(_2987_));
 sky130_fd_sc_hd__o211a_1 _6585_ (.A1(net66),
    .A2(_2987_),
    .B1(_2986_),
    .C1(net197),
    .X(_0048_));
 sky130_fd_sc_hd__and3_1 _6586_ (.A(\ann.X[25] ),
    .B(\ann.multiply_FF[25] ),
    .C(net196),
    .X(_2988_));
 sky130_fd_sc_hd__inv_2 _6587_ (.A(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__a21oi_1 _6588_ (.A1(\ann.multiply_FF[25] ),
    .A2(net196),
    .B1(\ann.X[25] ),
    .Y(_2990_));
 sky130_fd_sc_hd__a21o_1 _6589_ (.A1(\ann.multiply_FF[25] ),
    .A2(net196),
    .B1(\ann.X[25] ),
    .X(_2991_));
 sky130_fd_sc_hd__nor2_1 _6590_ (.A(_2988_),
    .B(_2990_),
    .Y(_2992_));
 sky130_fd_sc_hd__nor2_1 _6591_ (.A(_2977_),
    .B(_2981_),
    .Y(_2993_));
 sky130_fd_sc_hd__xnor2_1 _6592_ (.A(_2992_),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__and2_1 _6593_ (.A(\ann.bias[25] ),
    .B(\ann.sum[25] ),
    .X(_2995_));
 sky130_fd_sc_hd__or2_1 _6594_ (.A(\ann.bias[25] ),
    .B(\ann.sum[25] ),
    .X(_2996_));
 sky130_fd_sc_hd__and2b_1 _6595_ (.A_N(_2995_),
    .B(_2996_),
    .X(_2997_));
 sky130_fd_sc_hd__a21o_1 _6596_ (.A1(_2982_),
    .A2(_2985_),
    .B1(_2983_),
    .X(_2998_));
 sky130_fd_sc_hd__xnor2_1 _6597_ (.A(_2997_),
    .B(_2998_),
    .Y(_2999_));
 sky130_fd_sc_hd__nand2_1 _6598_ (.A(net62),
    .B(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__o211a_1 _6599_ (.A1(net62),
    .A2(_2994_),
    .B1(_3000_),
    .C1(net196),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _6600_ (.A1(\ann.multiply_FF[26] ),
    .A2(net196),
    .B1(\ann.X[26] ),
    .X(_3001_));
 sky130_fd_sc_hd__nand3_2 _6601_ (.A(\ann.X[26] ),
    .B(\ann.multiply_FF[26] ),
    .C(net196),
    .Y(_3002_));
 sky130_fd_sc_hd__nand2_1 _6602_ (.A(_3001_),
    .B(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__inv_2 _6603_ (.A(_3003_),
    .Y(_3004_));
 sky130_fd_sc_hd__o31a_1 _6604_ (.A1(_2977_),
    .A2(_2981_),
    .A3(_2988_),
    .B1(_2991_),
    .X(_3005_));
 sky130_fd_sc_hd__or2_1 _6605_ (.A(_3004_),
    .B(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__nand2_1 _6606_ (.A(_3004_),
    .B(_3005_),
    .Y(_3007_));
 sky130_fd_sc_hd__or2_1 _6607_ (.A(\ann.bias[26] ),
    .B(\ann.sum[26] ),
    .X(_3008_));
 sky130_fd_sc_hd__nand2_1 _6608_ (.A(\ann.bias[26] ),
    .B(\ann.sum[26] ),
    .Y(_3009_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(_3008_),
    .B(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__o21a_1 _6610_ (.A1(_2995_),
    .A2(_2998_),
    .B1(_2996_),
    .X(_3011_));
 sky130_fd_sc_hd__a21o_1 _6611_ (.A1(_3006_),
    .A2(_3007_),
    .B1(net62),
    .X(_3012_));
 sky130_fd_sc_hd__xnor2_1 _6612_ (.A(_3010_),
    .B(_3011_),
    .Y(_3013_));
 sky130_fd_sc_hd__o211a_1 _6613_ (.A1(net66),
    .A2(_3013_),
    .B1(_3012_),
    .C1(net196),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _6614_ (.A(\ann.bias[27] ),
    .B(\ann.sum[27] ),
    .X(_3014_));
 sky130_fd_sc_hd__nand2_1 _6615_ (.A(\ann.bias[27] ),
    .B(\ann.sum[27] ),
    .Y(_3015_));
 sky130_fd_sc_hd__inv_2 _6616_ (.A(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__nand2_1 _6617_ (.A(_3014_),
    .B(_3015_),
    .Y(_3017_));
 sky130_fd_sc_hd__a21boi_1 _6618_ (.A1(_3008_),
    .A2(_3011_),
    .B1_N(_3009_),
    .Y(_3018_));
 sky130_fd_sc_hd__xor2_1 _6619_ (.A(_3017_),
    .B(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__a21oi_1 _6620_ (.A1(\ann.multiply_FF[27] ),
    .A2(net196),
    .B1(\ann.X[27] ),
    .Y(_3020_));
 sky130_fd_sc_hd__and3_1 _6621_ (.A(\ann.X[27] ),
    .B(\ann.multiply_FF[27] ),
    .C(net196),
    .X(_3021_));
 sky130_fd_sc_hd__inv_2 _6622_ (.A(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__nor2_1 _6623_ (.A(_3020_),
    .B(_3021_),
    .Y(_3023_));
 sky130_fd_sc_hd__a21oi_1 _6624_ (.A1(_3002_),
    .A2(_3007_),
    .B1(_3023_),
    .Y(_3024_));
 sky130_fd_sc_hd__a31o_1 _6625_ (.A1(_3002_),
    .A2(_3007_),
    .A3(_3023_),
    .B1(net62),
    .X(_3025_));
 sky130_fd_sc_hd__or2_1 _6626_ (.A(_3024_),
    .B(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__o211a_1 _6627_ (.A1(net66),
    .A2(_3019_),
    .B1(_3026_),
    .C1(net196),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_1 _6628_ (.A(_3004_),
    .B(_3023_),
    .Y(_3027_));
 sky130_fd_sc_hd__and4_1 _6629_ (.A(_2979_),
    .B(_2992_),
    .C(_3004_),
    .D(_3023_),
    .X(_3028_));
 sky130_fd_sc_hd__o311ai_4 _6630_ (.A1(_2954_),
    .A2(_2956_),
    .A3(_2965_),
    .B1(_3028_),
    .C1(_2964_),
    .Y(_3029_));
 sky130_fd_sc_hd__a211o_1 _6631_ (.A1(_2976_),
    .A2(_2989_),
    .B1(_2990_),
    .C1(_3027_),
    .X(_3030_));
 sky130_fd_sc_hd__o211a_1 _6632_ (.A1(_3002_),
    .A2(_3020_),
    .B1(_3022_),
    .C1(_3030_),
    .X(_3031_));
 sky130_fd_sc_hd__a21oi_1 _6633_ (.A1(\ann.multiply_FF[28] ),
    .A2(net198),
    .B1(\ann.X[28] ),
    .Y(_3032_));
 sky130_fd_sc_hd__and3_1 _6634_ (.A(\ann.X[28] ),
    .B(\ann.multiply_FF[28] ),
    .C(net198),
    .X(_3033_));
 sky130_fd_sc_hd__or2_1 _6635_ (.A(_3032_),
    .B(_3033_),
    .X(_3034_));
 sky130_fd_sc_hd__and3_1 _6636_ (.A(_3029_),
    .B(_3031_),
    .C(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__a21oi_2 _6637_ (.A1(_3029_),
    .A2(_3031_),
    .B1(_3034_),
    .Y(_3036_));
 sky130_fd_sc_hd__or3_1 _6638_ (.A(net62),
    .B(_3035_),
    .C(_3036_),
    .X(_3037_));
 sky130_fd_sc_hd__nor2_1 _6639_ (.A(_3010_),
    .B(_3017_),
    .Y(_3038_));
 sky130_fd_sc_hd__and3_1 _6640_ (.A(_2985_),
    .B(_2997_),
    .C(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__or2_1 _6641_ (.A(_2983_),
    .B(_2995_),
    .X(_3040_));
 sky130_fd_sc_hd__a31o_1 _6642_ (.A1(\ann.bias[26] ),
    .A2(\ann.sum[26] ),
    .A3(_3014_),
    .B1(_3016_),
    .X(_3041_));
 sky130_fd_sc_hd__a31o_1 _6643_ (.A1(_2996_),
    .A2(_3038_),
    .A3(_3040_),
    .B1(_3041_),
    .X(_3042_));
 sky130_fd_sc_hd__a21oi_2 _6644_ (.A1(_2982_),
    .A2(_3039_),
    .B1(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__nor2_1 _6645_ (.A(\ann.bias[28] ),
    .B(\ann.sum[28] ),
    .Y(_3044_));
 sky130_fd_sc_hd__nand2_1 _6646_ (.A(\ann.bias[28] ),
    .B(\ann.sum[28] ),
    .Y(_3045_));
 sky130_fd_sc_hd__nand2b_1 _6647_ (.A_N(_3044_),
    .B(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__xor2_1 _6648_ (.A(_3043_),
    .B(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__nand2_1 _6649_ (.A(net62),
    .B(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__a21oi_1 _6650_ (.A1(_3037_),
    .A2(_3048_),
    .B1(net194),
    .Y(_0052_));
 sky130_fd_sc_hd__o21a_1 _6651_ (.A1(_3043_),
    .A2(_3044_),
    .B1(_3045_),
    .X(_3049_));
 sky130_fd_sc_hd__nor2_1 _6652_ (.A(\ann.bias[29] ),
    .B(\ann.sum[29] ),
    .Y(_3050_));
 sky130_fd_sc_hd__or2_1 _6653_ (.A(\ann.bias[29] ),
    .B(\ann.sum[29] ),
    .X(_3051_));
 sky130_fd_sc_hd__nand2_1 _6654_ (.A(\ann.bias[29] ),
    .B(\ann.sum[29] ),
    .Y(_3052_));
 sky130_fd_sc_hd__a21oi_1 _6655_ (.A1(_3051_),
    .A2(_3052_),
    .B1(_3049_),
    .Y(_3053_));
 sky130_fd_sc_hd__a31o_1 _6656_ (.A1(_3049_),
    .A2(_3051_),
    .A3(_3052_),
    .B1(net67),
    .X(_3054_));
 sky130_fd_sc_hd__a21oi_2 _6657_ (.A1(\ann.multiply_FF[29] ),
    .A2(net198),
    .B1(\ann.X[29] ),
    .Y(_3055_));
 sky130_fd_sc_hd__inv_2 _6658_ (.A(_3055_),
    .Y(_3056_));
 sky130_fd_sc_hd__and3_1 _6659_ (.A(\ann.X[29] ),
    .B(\ann.multiply_FF[29] ),
    .C(net198),
    .X(_3057_));
 sky130_fd_sc_hd__o22a_1 _6660_ (.A1(_3033_),
    .A2(_3036_),
    .B1(_3055_),
    .B2(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__nor4_1 _6661_ (.A(_3033_),
    .B(_3036_),
    .C(_3055_),
    .D(_3057_),
    .Y(_3059_));
 sky130_fd_sc_hd__o21a_1 _6662_ (.A1(_3053_),
    .A2(_3054_),
    .B1(net198),
    .X(_3060_));
 sky130_fd_sc_hd__o31a_1 _6663_ (.A1(net62),
    .A2(_3058_),
    .A3(_3059_),
    .B1(_3060_),
    .X(_0053_));
 sky130_fd_sc_hd__a21oi_1 _6664_ (.A1(\ann.multiply_FF[30] ),
    .A2(net199),
    .B1(\ann.X[30] ),
    .Y(_3061_));
 sky130_fd_sc_hd__and3_1 _6665_ (.A(\ann.X[30] ),
    .B(\ann.multiply_FF[30] ),
    .C(net199),
    .X(_3062_));
 sky130_fd_sc_hd__nor2_1 _6666_ (.A(_3061_),
    .B(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__or2_1 _6667_ (.A(_3033_),
    .B(_3057_),
    .X(_3064_));
 sky130_fd_sc_hd__o21a_1 _6668_ (.A1(_3036_),
    .A2(_3064_),
    .B1(_3056_),
    .X(_3065_));
 sky130_fd_sc_hd__nor2_1 _6669_ (.A(_3063_),
    .B(_3065_),
    .Y(_3066_));
 sky130_fd_sc_hd__o211a_1 _6670_ (.A1(_3036_),
    .A2(_3064_),
    .B1(_3063_),
    .C1(_3056_),
    .X(_3067_));
 sky130_fd_sc_hd__or3_1 _6671_ (.A(net62),
    .B(_3066_),
    .C(_3067_),
    .X(_3068_));
 sky130_fd_sc_hd__nand2_1 _6672_ (.A(\ann.bias[30] ),
    .B(\ann.sum[30] ),
    .Y(_3069_));
 sky130_fd_sc_hd__or2_1 _6673_ (.A(\ann.bias[30] ),
    .B(\ann.sum[30] ),
    .X(_3070_));
 sky130_fd_sc_hd__o21ai_2 _6674_ (.A1(_3049_),
    .A2(_3050_),
    .B1(_3052_),
    .Y(_3071_));
 sky130_fd_sc_hd__a21oi_1 _6675_ (.A1(_3069_),
    .A2(_3070_),
    .B1(_3071_),
    .Y(_3072_));
 sky130_fd_sc_hd__a31o_1 _6676_ (.A1(_3069_),
    .A2(_3070_),
    .A3(_3071_),
    .B1(net67),
    .X(_3073_));
 sky130_fd_sc_hd__or2_1 _6677_ (.A(_3072_),
    .B(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__a21oi_1 _6678_ (.A1(_3068_),
    .A2(_3074_),
    .B1(net194),
    .Y(_0055_));
 sky130_fd_sc_hd__a21bo_1 _6679_ (.A1(_3070_),
    .A2(_3071_),
    .B1_N(_3069_),
    .X(_3075_));
 sky130_fd_sc_hd__xnor2_1 _6680_ (.A(\ann.bias[31] ),
    .B(net59),
    .Y(_3076_));
 sky130_fd_sc_hd__xnor2_1 _6681_ (.A(_3075_),
    .B(_3076_),
    .Y(_3077_));
 sky130_fd_sc_hd__a21oi_1 _6682_ (.A1(\ann.multiply_FF[31] ),
    .A2(net198),
    .B1(\ann.X[31] ),
    .Y(_3078_));
 sky130_fd_sc_hd__and3_1 _6683_ (.A(\ann.X[31] ),
    .B(\ann.multiply_FF[31] ),
    .C(net198),
    .X(_3079_));
 sky130_fd_sc_hd__or4_1 _6684_ (.A(_3062_),
    .B(_3067_),
    .C(_3078_),
    .D(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__o22a_1 _6685_ (.A1(_3062_),
    .A2(_3067_),
    .B1(_3078_),
    .B2(_3079_),
    .X(_3081_));
 sky130_fd_sc_hd__or3b_1 _6686_ (.A(_3081_),
    .B(net62),
    .C_N(_3080_),
    .X(_3082_));
 sky130_fd_sc_hd__o211a_1 _6687_ (.A1(net67),
    .A2(_3077_),
    .B1(_3082_),
    .C1(net199),
    .X(_0056_));
 sky130_fd_sc_hd__o21ba_1 _6688_ (.A1(net402),
    .A2(net24),
    .B1_N(net789),
    .X(\ann.next_state[0] ));
 sky130_fd_sc_hd__a21o_1 _6689_ (.A1(_0565_),
    .A2(_0557_),
    .B1(_0558_),
    .X(\ann.next_state[1] ));
 sky130_fd_sc_hd__nor3_2 _6690_ (.A(net66),
    .B(net21),
    .C(net194),
    .Y(_0066_));
 sky130_fd_sc_hd__nor2_2 _6691_ (.A(net26),
    .B(net194),
    .Y(_0067_));
 sky130_fd_sc_hd__and2_1 _6692_ (.A(\ann.state[1] ),
    .B(\ann.state[0] ),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _6693_ (.A(\ann.multiply_out[0] ),
    .B(net201),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _6694_ (.A(\ann.multiply_out[1] ),
    .B(net202),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _6695_ (.A(\ann.multiply_out[2] ),
    .B(net202),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _6696_ (.A(\ann.multiply_out[3] ),
    .B(net204),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _6697_ (.A(\ann.multiply_out[4] ),
    .B(net205),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _6698_ (.A(\ann.multiply_out[5] ),
    .B(net208),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _6699_ (.A(\ann.multiply_out[6] ),
    .B(net208),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _6700_ (.A(\ann.multiply_out[7] ),
    .B(net208),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _6701_ (.A(\ann.multiply_out[8] ),
    .B(net208),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _6702_ (.A(\ann.multiply_out[9] ),
    .B(net208),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _6703_ (.A(\ann.multiply_out[10] ),
    .B(net208),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _6704_ (.A(\ann.multiply_out[11] ),
    .B(net208),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _6705_ (.A(\ann.multiply_out[12] ),
    .B(net207),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _6706_ (.A(\ann.multiply_out[13] ),
    .B(net207),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _6707_ (.A(\ann.multiply_out[14] ),
    .B(net207),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _6708_ (.A(\ann.multiply_out[15] ),
    .B(net207),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _6709_ (.A(\ann.multiply_out[16] ),
    .B(net202),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _6710_ (.A(\ann.multiply_out[17] ),
    .B(net202),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _6711_ (.A(\ann.multiply_out[18] ),
    .B(net199),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _6712_ (.A(\ann.multiply_out[19] ),
    .B(net200),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _6713_ (.A(\ann.multiply_out[20] ),
    .B(net200),
    .X(_0088_));
 sky130_fd_sc_hd__and2_1 _6714_ (.A(\ann.multiply_out[21] ),
    .B(net200),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _6715_ (.A(\ann.multiply_out[22] ),
    .B(net209),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _6716_ (.A(\ann.multiply_out[23] ),
    .B(net199),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _6717_ (.A(\ann.multiply_out[24] ),
    .B(net198),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _6718_ (.A(\ann.multiply_out[25] ),
    .B(net198),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _6719_ (.A(\ann.multiply_out[26] ),
    .B(net198),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _6720_ (.A(\ann.multiply_out[27] ),
    .B(net197),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _6721_ (.A(\ann.multiply_out[28] ),
    .B(net198),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _6722_ (.A(\ann.multiply_out[29] ),
    .B(net198),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _6723_ (.A(\ann.multiply_out[30] ),
    .B(net199),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _6724_ (.A(\ann.multiply_out[31] ),
    .B(net199),
    .X(_0099_));
 sky130_fd_sc_hd__o22a_1 _6725_ (.A1(net103),
    .A2(\ann.ReLU_out[9][15] ),
    .B1(\ann.ReLU_out[9][14] ),
    .B2(net102),
    .X(_3083_));
 sky130_fd_sc_hd__a22o_1 _6726_ (.A1(net102),
    .A2(\ann.ReLU_out[9][14] ),
    .B1(\ann.ReLU_out[9][13] ),
    .B2(net101),
    .X(_3084_));
 sky130_fd_sc_hd__a22o_1 _6727_ (.A1(\ann.temp[11] ),
    .A2(_0704_),
    .B1(_0705_),
    .B2(\ann.temp[10] ),
    .X(_3085_));
 sky130_fd_sc_hd__a22o_1 _6728_ (.A1(\ann.temp[9] ),
    .A2(_0706_),
    .B1(_0707_),
    .B2(net189),
    .X(_3086_));
 sky130_fd_sc_hd__o22a_1 _6729_ (.A1(\ann.temp[10] ),
    .A2(_0705_),
    .B1(_0706_),
    .B2(\ann.temp[9] ),
    .X(_3087_));
 sky130_fd_sc_hd__a21oi_1 _6730_ (.A1(_3086_),
    .A2(_3087_),
    .B1(_3085_),
    .Y(_3088_));
 sky130_fd_sc_hd__nor2_1 _6731_ (.A(\ann.temp[11] ),
    .B(_0704_),
    .Y(_3089_));
 sky130_fd_sc_hd__and2_1 _6732_ (.A(net100),
    .B(\ann.ReLU_out[9][12] ),
    .X(_3090_));
 sky130_fd_sc_hd__or3_1 _6733_ (.A(_3088_),
    .B(_3089_),
    .C(_3090_),
    .X(_3091_));
 sky130_fd_sc_hd__o221a_1 _6734_ (.A1(net101),
    .A2(\ann.ReLU_out[9][13] ),
    .B1(\ann.ReLU_out[9][12] ),
    .B2(net100),
    .C1(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__or2_1 _6735_ (.A(_3084_),
    .B(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__a22o_1 _6736_ (.A1(net103),
    .A2(\ann.ReLU_out[9][15] ),
    .B1(_3083_),
    .B2(_3093_),
    .X(_3094_));
 sky130_fd_sc_hd__or2_1 _6737_ (.A(net98),
    .B(\ann.ReLU_out[9][6] ),
    .X(_3095_));
 sky130_fd_sc_hd__or2_1 _6738_ (.A(net93),
    .B(\ann.ReLU_out[9][1] ),
    .X(_3096_));
 sky130_fd_sc_hd__a22o_1 _6739_ (.A1(net94),
    .A2(\ann.ReLU_out[9][2] ),
    .B1(\ann.ReLU_out[9][1] ),
    .B2(net93),
    .X(_3097_));
 sky130_fd_sc_hd__a31o_1 _6740_ (.A1(_0661_),
    .A2(\ann.ReLU_out[9][0] ),
    .A3(_3096_),
    .B1(_3097_),
    .X(_3098_));
 sky130_fd_sc_hd__o221a_1 _6741_ (.A1(net95),
    .A2(\ann.ReLU_out[9][3] ),
    .B1(net577),
    .B2(net94),
    .C1(_3098_),
    .X(_3099_));
 sky130_fd_sc_hd__a221o_1 _6742_ (.A1(net96),
    .A2(net606),
    .B1(\ann.ReLU_out[9][3] ),
    .B2(net95),
    .C1(_3099_),
    .X(_3100_));
 sky130_fd_sc_hd__o221a_1 _6743_ (.A1(net97),
    .A2(\ann.ReLU_out[9][5] ),
    .B1(net606),
    .B2(net96),
    .C1(_3100_),
    .X(_3101_));
 sky130_fd_sc_hd__a221o_1 _6744_ (.A1(net98),
    .A2(\ann.ReLU_out[9][6] ),
    .B1(\ann.ReLU_out[9][5] ),
    .B2(net97),
    .C1(_3101_),
    .X(_3102_));
 sky130_fd_sc_hd__a22o_1 _6745_ (.A1(net99),
    .A2(\ann.ReLU_out[9][7] ),
    .B1(_3095_),
    .B2(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__o21a_2 _6746_ (.A1(net99),
    .A2(\ann.ReLU_out[9][7] ),
    .B1(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__o221a_1 _6747_ (.A1(\ann.temp[15] ),
    .A2(_0703_),
    .B1(_0707_),
    .B2(net189),
    .C1(_3083_),
    .X(_3105_));
 sky130_fd_sc_hd__or2_1 _6748_ (.A(_3084_),
    .B(_3090_),
    .X(_3106_));
 sky130_fd_sc_hd__or4b_1 _6749_ (.A(_3086_),
    .B(_3089_),
    .C(_3106_),
    .D_N(_3087_),
    .X(_3107_));
 sky130_fd_sc_hd__o221a_1 _6750_ (.A1(net101),
    .A2(\ann.ReLU_out[9][13] ),
    .B1(\ann.ReLU_out[9][12] ),
    .B2(net100),
    .C1(_3105_),
    .X(_3108_));
 sky130_fd_sc_hd__or4b_1 _6751_ (.A(_3085_),
    .B(_3104_),
    .C(_3107_),
    .D_N(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__nand2_1 _6752_ (.A(_3094_),
    .B(_3109_),
    .Y(_3110_));
 sky130_fd_sc_hd__a22o_1 _6753_ (.A1(net188),
    .A2(_0701_),
    .B1(_0702_),
    .B2(\ann.temp[16] ),
    .X(_3111_));
 sky130_fd_sc_hd__o22a_1 _6754_ (.A1(net187),
    .A2(_0700_),
    .B1(_0701_),
    .B2(net188),
    .X(_3112_));
 sky130_fd_sc_hd__xnor2_1 _6755_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[9][19] ),
    .Y(_3113_));
 sky130_fd_sc_hd__o221a_1 _6756_ (.A1(_0640_),
    .A2(\ann.ReLU_out[9][18] ),
    .B1(_0702_),
    .B2(\ann.temp[16] ),
    .C1(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__and4b_1 _6757_ (.A_N(_3111_),
    .B(_3112_),
    .C(_3114_),
    .D(_3110_),
    .X(_3115_));
 sky130_fd_sc_hd__a2bb2o_1 _6758_ (.A1_N(\ann.ReLU_out[9][25] ),
    .A2_N(_0574_),
    .B1(net184),
    .B2(_0575_),
    .X(_3116_));
 sky130_fd_sc_hd__a22o_1 _6759_ (.A1(\ann.ReLU_out[9][26] ),
    .A2(_0573_),
    .B1(\ann.ReLU_out[9][25] ),
    .B2(_0574_),
    .X(_3117_));
 sky130_fd_sc_hd__o22a_1 _6760_ (.A1(net184),
    .A2(_0575_),
    .B1(_0576_),
    .B2(net185),
    .X(_3118_));
 sky130_fd_sc_hd__inv_2 _6761_ (.A(_3118_),
    .Y(_3119_));
 sky130_fd_sc_hd__a221o_1 _6762_ (.A1(_0576_),
    .A2(net185),
    .B1(_0577_),
    .B2(net186),
    .C1(_3119_),
    .X(_3120_));
 sky130_fd_sc_hd__a2bb2o_1 _6763_ (.A1_N(\ann.ReLU_out[9][29] ),
    .A2_N(_0569_),
    .B1(_0570_),
    .B2(\ann.temp[28] ),
    .X(_3121_));
 sky130_fd_sc_hd__nand2_1 _6764_ (.A(\ann.ReLU_out[9][29] ),
    .B(_0569_),
    .Y(_3122_));
 sky130_fd_sc_hd__nor2_1 _6765_ (.A(_0570_),
    .B(\ann.temp[28] ),
    .Y(_3123_));
 sky130_fd_sc_hd__or3b_1 _6766_ (.A(_3123_),
    .B(_3121_),
    .C_N(_3122_),
    .X(_3124_));
 sky130_fd_sc_hd__or2_1 _6767_ (.A(\ann.ReLU_out[9][21] ),
    .B(_0579_),
    .X(_3125_));
 sky130_fd_sc_hd__a22o_1 _6768_ (.A1(\ann.ReLU_out[9][21] ),
    .A2(_0579_),
    .B1(_0580_),
    .B2(\ann.ReLU_out[9][20] ),
    .X(_3126_));
 sky130_fd_sc_hd__o22ai_1 _6769_ (.A1(_0580_),
    .A2(\ann.ReLU_out[9][20] ),
    .B1(_0639_),
    .B2(\ann.ReLU_out[9][19] ),
    .Y(_3127_));
 sky130_fd_sc_hd__nor2_1 _6770_ (.A(net104),
    .B(\ann.ReLU_out[9][30] ),
    .Y(_3128_));
 sky130_fd_sc_hd__o22ai_2 _6771_ (.A1(\ann.ReLU_out[9][27] ),
    .A2(_0572_),
    .B1(\ann.ReLU_out[9][26] ),
    .B2(_0573_),
    .Y(_3129_));
 sky130_fd_sc_hd__a221o_1 _6772_ (.A1(net104),
    .A2(\ann.ReLU_out[9][30] ),
    .B1(\ann.ReLU_out[9][27] ),
    .B2(_0572_),
    .C1(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__a2111o_1 _6773_ (.A1(\ann.ReLU_out[9][22] ),
    .A2(_0578_),
    .B1(_3127_),
    .C1(_3128_),
    .D1(_3130_),
    .X(_3131_));
 sky130_fd_sc_hd__or4b_1 _6774_ (.A(_3124_),
    .B(_3126_),
    .C(_3131_),
    .D_N(_3125_),
    .X(_3132_));
 sky130_fd_sc_hd__or4_2 _6775_ (.A(_3116_),
    .B(_3117_),
    .C(_3120_),
    .D(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__a22o_1 _6776_ (.A1(net187),
    .A2(_0700_),
    .B1(_3111_),
    .B2(_3112_),
    .X(_3134_));
 sky130_fd_sc_hd__a211o_1 _6777_ (.A1(_3113_),
    .A2(_3134_),
    .B1(_3133_),
    .C1(_3115_),
    .X(_3135_));
 sky130_fd_sc_hd__o2bb2a_1 _6778_ (.A1_N(_3125_),
    .A2_N(_3126_),
    .B1(_0577_),
    .B2(net186),
    .X(_3136_));
 sky130_fd_sc_hd__a221o_1 _6779_ (.A1(_0576_),
    .A2(net185),
    .B1(_0577_),
    .B2(net186),
    .C1(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__a21oi_1 _6780_ (.A1(_3118_),
    .A2(_3137_),
    .B1(_3116_),
    .Y(_3138_));
 sky130_fd_sc_hd__o21bai_1 _6781_ (.A1(_3117_),
    .A2(_3138_),
    .B1_N(_3129_),
    .Y(_3139_));
 sky130_fd_sc_hd__a21oi_1 _6782_ (.A1(\ann.ReLU_out[9][27] ),
    .A2(_0572_),
    .B1(_3124_),
    .Y(_3140_));
 sky130_fd_sc_hd__a221o_1 _6783_ (.A1(_3121_),
    .A2(_3122_),
    .B1(_3139_),
    .B2(_3140_),
    .C1(_3128_),
    .X(_3141_));
 sky130_fd_sc_hd__o211a_4 _6784_ (.A1(net788),
    .A2(_0568_),
    .B1(_3135_),
    .C1(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__o22a_1 _6785_ (.A1(net103),
    .A2(\ann.ReLU_out[8][15] ),
    .B1(\ann.ReLU_out[8][14] ),
    .B2(net102),
    .X(_3143_));
 sky130_fd_sc_hd__a22o_1 _6786_ (.A1(net102),
    .A2(\ann.ReLU_out[8][14] ),
    .B1(\ann.ReLU_out[8][13] ),
    .B2(net101),
    .X(_3144_));
 sky130_fd_sc_hd__o22a_1 _6787_ (.A1(net101),
    .A2(\ann.ReLU_out[8][13] ),
    .B1(\ann.ReLU_out[8][12] ),
    .B2(net100),
    .X(_3145_));
 sky130_fd_sc_hd__a22o_1 _6788_ (.A1(\ann.temp[11] ),
    .A2(_0696_),
    .B1(_0697_),
    .B2(\ann.temp[10] ),
    .X(_3146_));
 sky130_fd_sc_hd__a22o_1 _6789_ (.A1(\ann.temp[9] ),
    .A2(_0698_),
    .B1(_0699_),
    .B2(net189),
    .X(_3147_));
 sky130_fd_sc_hd__o22a_1 _6790_ (.A1(\ann.temp[10] ),
    .A2(_0697_),
    .B1(_0698_),
    .B2(\ann.temp[9] ),
    .X(_3148_));
 sky130_fd_sc_hd__a21oi_1 _6791_ (.A1(_3147_),
    .A2(_3148_),
    .B1(_3146_),
    .Y(_3149_));
 sky130_fd_sc_hd__nor2_1 _6792_ (.A(\ann.temp[11] ),
    .B(_0696_),
    .Y(_3150_));
 sky130_fd_sc_hd__and2_1 _6793_ (.A(net100),
    .B(\ann.ReLU_out[8][12] ),
    .X(_3151_));
 sky130_fd_sc_hd__o31a_1 _6794_ (.A1(_3149_),
    .A2(_3150_),
    .A3(_3151_),
    .B1(_3145_),
    .X(_3152_));
 sky130_fd_sc_hd__or2_1 _6795_ (.A(_3144_),
    .B(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__a22o_1 _6796_ (.A1(net103),
    .A2(\ann.ReLU_out[8][15] ),
    .B1(_3143_),
    .B2(_3153_),
    .X(_3154_));
 sky130_fd_sc_hd__or2_1 _6797_ (.A(net98),
    .B(\ann.ReLU_out[8][6] ),
    .X(_3155_));
 sky130_fd_sc_hd__or2_1 _6798_ (.A(net93),
    .B(\ann.ReLU_out[8][1] ),
    .X(_3156_));
 sky130_fd_sc_hd__a22o_1 _6799_ (.A1(net94),
    .A2(\ann.ReLU_out[8][2] ),
    .B1(\ann.ReLU_out[8][1] ),
    .B2(net93),
    .X(_3157_));
 sky130_fd_sc_hd__a31o_1 _6800_ (.A1(_0661_),
    .A2(\ann.ReLU_out[8][0] ),
    .A3(_3156_),
    .B1(_3157_),
    .X(_3158_));
 sky130_fd_sc_hd__o221a_1 _6801_ (.A1(net95),
    .A2(\ann.ReLU_out[8][3] ),
    .B1(\ann.ReLU_out[8][2] ),
    .B2(net94),
    .C1(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__a221o_1 _6802_ (.A1(net96),
    .A2(\ann.ReLU_out[8][4] ),
    .B1(\ann.ReLU_out[8][3] ),
    .B2(net95),
    .C1(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__o221a_1 _6803_ (.A1(net97),
    .A2(\ann.ReLU_out[8][5] ),
    .B1(\ann.ReLU_out[8][4] ),
    .B2(net96),
    .C1(_3160_),
    .X(_3161_));
 sky130_fd_sc_hd__a221o_1 _6804_ (.A1(net98),
    .A2(\ann.ReLU_out[8][6] ),
    .B1(\ann.ReLU_out[8][5] ),
    .B2(net97),
    .C1(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__a22o_1 _6805_ (.A1(net99),
    .A2(\ann.ReLU_out[8][7] ),
    .B1(_3155_),
    .B2(_3162_),
    .X(_3163_));
 sky130_fd_sc_hd__o21a_1 _6806_ (.A1(net99),
    .A2(\ann.ReLU_out[8][7] ),
    .B1(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__o221a_1 _6807_ (.A1(\ann.temp[15] ),
    .A2(_0695_),
    .B1(_0699_),
    .B2(net189),
    .C1(_3143_),
    .X(_3165_));
 sky130_fd_sc_hd__or2_1 _6808_ (.A(_3144_),
    .B(_3151_),
    .X(_3166_));
 sky130_fd_sc_hd__or4b_1 _6809_ (.A(_3147_),
    .B(_3150_),
    .C(_3166_),
    .D_N(_3148_),
    .X(_3167_));
 sky130_fd_sc_hd__nand2_1 _6810_ (.A(_3145_),
    .B(_3165_),
    .Y(_3168_));
 sky130_fd_sc_hd__o41a_1 _6811_ (.A1(_3146_),
    .A2(_3164_),
    .A3(_3167_),
    .A4(_3168_),
    .B1(_3154_),
    .X(_3169_));
 sky130_fd_sc_hd__a2bb2o_1 _6812_ (.A1_N(\ann.ReLU_out[8][16] ),
    .A2_N(_0643_),
    .B1(net188),
    .B2(_0694_),
    .X(_3170_));
 sky130_fd_sc_hd__nor2_1 _6813_ (.A(_0640_),
    .B(\ann.ReLU_out[8][18] ),
    .Y(_3171_));
 sky130_fd_sc_hd__xor2_1 _6814_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[8][19] ),
    .X(_3172_));
 sky130_fd_sc_hd__a221o_1 _6815_ (.A1(_0640_),
    .A2(\ann.ReLU_out[8][18] ),
    .B1(\ann.ReLU_out[8][17] ),
    .B2(_0642_),
    .C1(_3170_),
    .X(_3173_));
 sky130_fd_sc_hd__a211o_1 _6816_ (.A1(_0643_),
    .A2(\ann.ReLU_out[8][16] ),
    .B1(_3171_),
    .C1(_3172_),
    .X(_3174_));
 sky130_fd_sc_hd__nor3_1 _6817_ (.A(_3169_),
    .B(_3173_),
    .C(_3174_),
    .Y(_3175_));
 sky130_fd_sc_hd__o221a_1 _6818_ (.A1(net187),
    .A2(_0693_),
    .B1(_0694_),
    .B2(net188),
    .C1(_3170_),
    .X(_3176_));
 sky130_fd_sc_hd__o21ba_1 _6819_ (.A1(_3171_),
    .A2(_3176_),
    .B1_N(_3172_),
    .X(_3177_));
 sky130_fd_sc_hd__o22a_1 _6820_ (.A1(net184),
    .A2(_0584_),
    .B1(_0585_),
    .B2(net185),
    .X(_3178_));
 sky130_fd_sc_hd__inv_2 _6821_ (.A(_3178_),
    .Y(_3179_));
 sky130_fd_sc_hd__a221o_1 _6822_ (.A1(net185),
    .A2(_0585_),
    .B1(_0586_),
    .B2(net186),
    .C1(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__a22o_1 _6823_ (.A1(net183),
    .A2(_0583_),
    .B1(_0584_),
    .B2(net184),
    .X(_3181_));
 sky130_fd_sc_hd__a22o_1 _6824_ (.A1(_0571_),
    .A2(\ann.ReLU_out[8][28] ),
    .B1(\ann.ReLU_out[8][27] ),
    .B2(_0572_),
    .X(_3182_));
 sky130_fd_sc_hd__a2bb2o_1 _6825_ (.A1_N(_0572_),
    .A2_N(\ann.ReLU_out[8][27] ),
    .B1(_0582_),
    .B2(net182),
    .X(_3183_));
 sky130_fd_sc_hd__o22a_1 _6826_ (.A1(net182),
    .A2(_0582_),
    .B1(_0583_),
    .B2(net183),
    .X(_3184_));
 sky130_fd_sc_hd__inv_2 _6827_ (.A(_3184_),
    .Y(_3185_));
 sky130_fd_sc_hd__a22o_1 _6828_ (.A1(_0579_),
    .A2(\ann.ReLU_out[8][21] ),
    .B1(\ann.ReLU_out[8][20] ),
    .B2(_0580_),
    .X(_3186_));
 sky130_fd_sc_hd__a2bb2o_1 _6829_ (.A1_N(\ann.ReLU_out[8][28] ),
    .A2_N(_0571_),
    .B1(\ann.temp[29] ),
    .B2(_0581_),
    .X(_3187_));
 sky130_fd_sc_hd__or4_1 _6830_ (.A(_3183_),
    .B(_3185_),
    .C(_3186_),
    .D(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__nor2_1 _6831_ (.A(net186),
    .B(_0586_),
    .Y(_3189_));
 sky130_fd_sc_hd__nand2_1 _6832_ (.A(\ann.temp[21] ),
    .B(_0587_),
    .Y(_3190_));
 sky130_fd_sc_hd__nand2_1 _6833_ (.A(net104),
    .B(net610),
    .Y(_3191_));
 sky130_fd_sc_hd__o21ai_1 _6834_ (.A1(_0639_),
    .A2(\ann.ReLU_out[8][19] ),
    .B1(_3191_),
    .Y(_3192_));
 sky130_fd_sc_hd__nor2_1 _6835_ (.A(net104),
    .B(\ann.ReLU_out[8][30] ),
    .Y(_3193_));
 sky130_fd_sc_hd__a221o_1 _6836_ (.A1(_0569_),
    .A2(\ann.ReLU_out[8][29] ),
    .B1(_0588_),
    .B2(\ann.temp[20] ),
    .C1(_3182_),
    .X(_3194_));
 sky130_fd_sc_hd__a2111o_1 _6837_ (.A1(\ann.temp[21] ),
    .A2(_0587_),
    .B1(_3189_),
    .C1(_3193_),
    .D1(_3194_),
    .X(_3195_));
 sky130_fd_sc_hd__or4_1 _6838_ (.A(_3180_),
    .B(_3181_),
    .C(_3192_),
    .D(_3195_),
    .X(_3196_));
 sky130_fd_sc_hd__or4_1 _6839_ (.A(_3175_),
    .B(_3177_),
    .C(_3188_),
    .D(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__a21oi_1 _6840_ (.A1(_3186_),
    .A2(_3190_),
    .B1(_3189_),
    .Y(_3198_));
 sky130_fd_sc_hd__a221o_1 _6841_ (.A1(net185),
    .A2(_0585_),
    .B1(_0586_),
    .B2(net186),
    .C1(_3198_),
    .X(_3199_));
 sky130_fd_sc_hd__a21o_1 _6842_ (.A1(_3178_),
    .A2(_3199_),
    .B1(_3181_),
    .X(_3200_));
 sky130_fd_sc_hd__a21oi_1 _6843_ (.A1(_3184_),
    .A2(_3200_),
    .B1(_3183_),
    .Y(_3201_));
 sky130_fd_sc_hd__nor2_1 _6844_ (.A(_3182_),
    .B(_3201_),
    .Y(_3202_));
 sky130_fd_sc_hd__o22a_1 _6845_ (.A1(\ann.temp[29] ),
    .A2(_0581_),
    .B1(_3187_),
    .B2(_3202_),
    .X(_3203_));
 sky130_fd_sc_hd__o211a_1 _6846_ (.A1(_3193_),
    .A2(_3203_),
    .B1(_3197_),
    .C1(_3191_),
    .X(_3204_));
 sky130_fd_sc_hd__o22a_1 _6847_ (.A1(net103),
    .A2(\ann.ReLU_out[7][15] ),
    .B1(\ann.ReLU_out[7][14] ),
    .B2(net102),
    .X(_3205_));
 sky130_fd_sc_hd__a22o_1 _6848_ (.A1(net102),
    .A2(\ann.ReLU_out[7][14] ),
    .B1(\ann.ReLU_out[7][13] ),
    .B2(net101),
    .X(_3206_));
 sky130_fd_sc_hd__o22a_1 _6849_ (.A1(net101),
    .A2(\ann.ReLU_out[7][13] ),
    .B1(\ann.ReLU_out[7][12] ),
    .B2(net100),
    .X(_3207_));
 sky130_fd_sc_hd__a22o_1 _6850_ (.A1(\ann.temp[11] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\ann.temp[10] ),
    .X(_3208_));
 sky130_fd_sc_hd__a22o_1 _6851_ (.A1(\ann.temp[9] ),
    .A2(_0691_),
    .B1(_0692_),
    .B2(net189),
    .X(_3209_));
 sky130_fd_sc_hd__o22a_1 _6852_ (.A1(\ann.temp[10] ),
    .A2(_0690_),
    .B1(_0691_),
    .B2(\ann.temp[9] ),
    .X(_3210_));
 sky130_fd_sc_hd__a21oi_1 _6853_ (.A1(_3209_),
    .A2(_3210_),
    .B1(_3208_),
    .Y(_3211_));
 sky130_fd_sc_hd__nor2_1 _6854_ (.A(\ann.temp[11] ),
    .B(_0689_),
    .Y(_3212_));
 sky130_fd_sc_hd__and2_1 _6855_ (.A(net100),
    .B(\ann.ReLU_out[7][12] ),
    .X(_3213_));
 sky130_fd_sc_hd__o31a_1 _6856_ (.A1(_3211_),
    .A2(_3212_),
    .A3(_3213_),
    .B1(_3207_),
    .X(_3214_));
 sky130_fd_sc_hd__or2_1 _6857_ (.A(_3206_),
    .B(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__a22o_1 _6858_ (.A1(net103),
    .A2(\ann.ReLU_out[7][15] ),
    .B1(_3205_),
    .B2(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__or2_1 _6859_ (.A(net98),
    .B(\ann.ReLU_out[7][6] ),
    .X(_3217_));
 sky130_fd_sc_hd__or2_1 _6860_ (.A(net93),
    .B(\ann.ReLU_out[7][1] ),
    .X(_3218_));
 sky130_fd_sc_hd__a22o_1 _6861_ (.A1(net94),
    .A2(\ann.ReLU_out[7][2] ),
    .B1(\ann.ReLU_out[7][1] ),
    .B2(net93),
    .X(_3219_));
 sky130_fd_sc_hd__a31o_1 _6862_ (.A1(_0661_),
    .A2(\ann.ReLU_out[7][0] ),
    .A3(_3218_),
    .B1(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__o221a_1 _6863_ (.A1(net95),
    .A2(\ann.ReLU_out[7][3] ),
    .B1(\ann.ReLU_out[7][2] ),
    .B2(net94),
    .C1(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__a221o_1 _6864_ (.A1(net96),
    .A2(\ann.ReLU_out[7][4] ),
    .B1(\ann.ReLU_out[7][3] ),
    .B2(net95),
    .C1(_3221_),
    .X(_3222_));
 sky130_fd_sc_hd__o221a_1 _6865_ (.A1(net97),
    .A2(\ann.ReLU_out[7][5] ),
    .B1(\ann.ReLU_out[7][4] ),
    .B2(net96),
    .C1(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__a221o_1 _6866_ (.A1(net98),
    .A2(\ann.ReLU_out[7][6] ),
    .B1(\ann.ReLU_out[7][5] ),
    .B2(net97),
    .C1(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__a22o_1 _6867_ (.A1(net99),
    .A2(\ann.ReLU_out[7][7] ),
    .B1(_3217_),
    .B2(_3224_),
    .X(_3225_));
 sky130_fd_sc_hd__o21a_1 _6868_ (.A1(net99),
    .A2(\ann.ReLU_out[7][7] ),
    .B1(_3225_),
    .X(_3226_));
 sky130_fd_sc_hd__o221a_1 _6869_ (.A1(\ann.temp[15] ),
    .A2(_0688_),
    .B1(_0692_),
    .B2(net189),
    .C1(_3205_),
    .X(_3227_));
 sky130_fd_sc_hd__or2_1 _6870_ (.A(_3206_),
    .B(_3213_),
    .X(_3228_));
 sky130_fd_sc_hd__or4b_1 _6871_ (.A(_3209_),
    .B(_3212_),
    .C(_3228_),
    .D_N(_3210_),
    .X(_3229_));
 sky130_fd_sc_hd__nand2_1 _6872_ (.A(_3207_),
    .B(_3227_),
    .Y(_3230_));
 sky130_fd_sc_hd__o41a_1 _6873_ (.A1(_3208_),
    .A2(_3226_),
    .A3(_3229_),
    .A4(_3230_),
    .B1(_3216_),
    .X(_3231_));
 sky130_fd_sc_hd__a2bb2o_1 _6874_ (.A1_N(\ann.ReLU_out[7][16] ),
    .A2_N(_0643_),
    .B1(net188),
    .B2(_0687_),
    .X(_3232_));
 sky130_fd_sc_hd__nor2_1 _6875_ (.A(_0640_),
    .B(\ann.ReLU_out[7][18] ),
    .Y(_3233_));
 sky130_fd_sc_hd__xor2_1 _6876_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[7][19] ),
    .X(_3234_));
 sky130_fd_sc_hd__a221o_1 _6877_ (.A1(_0640_),
    .A2(\ann.ReLU_out[7][18] ),
    .B1(\ann.ReLU_out[7][17] ),
    .B2(_0642_),
    .C1(_3232_),
    .X(_3235_));
 sky130_fd_sc_hd__a211o_1 _6878_ (.A1(_0643_),
    .A2(\ann.ReLU_out[7][16] ),
    .B1(_3233_),
    .C1(_3234_),
    .X(_3236_));
 sky130_fd_sc_hd__nor3_1 _6879_ (.A(_3231_),
    .B(_3235_),
    .C(_3236_),
    .Y(_3237_));
 sky130_fd_sc_hd__o221a_1 _6880_ (.A1(net187),
    .A2(_0686_),
    .B1(_0687_),
    .B2(net188),
    .C1(_3232_),
    .X(_3238_));
 sky130_fd_sc_hd__o21ba_1 _6881_ (.A1(_3233_),
    .A2(_3238_),
    .B1_N(_3234_),
    .X(_3239_));
 sky130_fd_sc_hd__o22a_1 _6882_ (.A1(net184),
    .A2(_0592_),
    .B1(_0593_),
    .B2(net185),
    .X(_3240_));
 sky130_fd_sc_hd__inv_2 _6883_ (.A(_3240_),
    .Y(_3241_));
 sky130_fd_sc_hd__a221o_1 _6884_ (.A1(net185),
    .A2(_0593_),
    .B1(_0594_),
    .B2(net186),
    .C1(_3241_),
    .X(_3242_));
 sky130_fd_sc_hd__a22o_1 _6885_ (.A1(net183),
    .A2(_0591_),
    .B1(_0592_),
    .B2(net184),
    .X(_3243_));
 sky130_fd_sc_hd__a22o_1 _6886_ (.A1(_0571_),
    .A2(\ann.ReLU_out[7][28] ),
    .B1(\ann.ReLU_out[7][27] ),
    .B2(_0572_),
    .X(_3244_));
 sky130_fd_sc_hd__a2bb2o_1 _6887_ (.A1_N(_0572_),
    .A2_N(\ann.ReLU_out[7][27] ),
    .B1(_0590_),
    .B2(net182),
    .X(_3245_));
 sky130_fd_sc_hd__o22a_1 _6888_ (.A1(net182),
    .A2(_0590_),
    .B1(_0591_),
    .B2(net183),
    .X(_3246_));
 sky130_fd_sc_hd__inv_2 _6889_ (.A(_3246_),
    .Y(_3247_));
 sky130_fd_sc_hd__a22o_1 _6890_ (.A1(_0579_),
    .A2(\ann.ReLU_out[7][21] ),
    .B1(\ann.ReLU_out[7][20] ),
    .B2(_0580_),
    .X(_3248_));
 sky130_fd_sc_hd__a2bb2o_1 _6891_ (.A1_N(\ann.ReLU_out[7][28] ),
    .A2_N(_0571_),
    .B1(\ann.temp[29] ),
    .B2(_0589_),
    .X(_3249_));
 sky130_fd_sc_hd__or4_1 _6892_ (.A(_3245_),
    .B(_3247_),
    .C(_3248_),
    .D(_3249_),
    .X(_3250_));
 sky130_fd_sc_hd__nor2_1 _6893_ (.A(net186),
    .B(_0594_),
    .Y(_3251_));
 sky130_fd_sc_hd__nand2_1 _6894_ (.A(\ann.temp[21] ),
    .B(_0595_),
    .Y(_3252_));
 sky130_fd_sc_hd__nand2_1 _6895_ (.A(net104),
    .B(\ann.ReLU_out[7][30] ),
    .Y(_3253_));
 sky130_fd_sc_hd__o21ai_1 _6896_ (.A1(_0639_),
    .A2(\ann.ReLU_out[7][19] ),
    .B1(_3253_),
    .Y(_3254_));
 sky130_fd_sc_hd__nor2_1 _6897_ (.A(net104),
    .B(\ann.ReLU_out[7][30] ),
    .Y(_3255_));
 sky130_fd_sc_hd__a221o_1 _6898_ (.A1(_0569_),
    .A2(\ann.ReLU_out[7][29] ),
    .B1(_0596_),
    .B2(\ann.temp[20] ),
    .C1(_3244_),
    .X(_3256_));
 sky130_fd_sc_hd__a2111o_1 _6899_ (.A1(\ann.temp[21] ),
    .A2(_0595_),
    .B1(_3251_),
    .C1(_3255_),
    .D1(_3256_),
    .X(_3257_));
 sky130_fd_sc_hd__or4_1 _6900_ (.A(_3242_),
    .B(_3243_),
    .C(_3254_),
    .D(_3257_),
    .X(_3258_));
 sky130_fd_sc_hd__or4_1 _6901_ (.A(_3237_),
    .B(_3239_),
    .C(_3250_),
    .D(_3258_),
    .X(_3259_));
 sky130_fd_sc_hd__a21oi_1 _6902_ (.A1(_3248_),
    .A2(_3252_),
    .B1(_3251_),
    .Y(_3260_));
 sky130_fd_sc_hd__a221o_1 _6903_ (.A1(net185),
    .A2(_0593_),
    .B1(_0594_),
    .B2(net186),
    .C1(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__a21o_1 _6904_ (.A1(_3240_),
    .A2(_3261_),
    .B1(_3243_),
    .X(_3262_));
 sky130_fd_sc_hd__a21oi_1 _6905_ (.A1(_3246_),
    .A2(_3262_),
    .B1(_3245_),
    .Y(_3263_));
 sky130_fd_sc_hd__nor2_1 _6906_ (.A(_3244_),
    .B(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__o22a_1 _6907_ (.A1(\ann.temp[29] ),
    .A2(_0589_),
    .B1(_3249_),
    .B2(_3264_),
    .X(_3265_));
 sky130_fd_sc_hd__o211ai_1 _6908_ (.A1(_3255_),
    .A2(_3265_),
    .B1(_3259_),
    .C1(_3253_),
    .Y(_3266_));
 sky130_fd_sc_hd__nor2_1 _6909_ (.A(\ann.temp[30] ),
    .B(_0597_),
    .Y(_3267_));
 sky130_fd_sc_hd__a22o_1 _6910_ (.A1(\ann.temp[27] ),
    .A2(_0598_),
    .B1(_0599_),
    .B2(net182),
    .X(_3268_));
 sky130_fd_sc_hd__o22a_1 _6911_ (.A1(net182),
    .A2(_0599_),
    .B1(_0600_),
    .B2(net183),
    .X(_3269_));
 sky130_fd_sc_hd__a22o_1 _6912_ (.A1(net183),
    .A2(_0600_),
    .B1(_0601_),
    .B2(net184),
    .X(_3270_));
 sky130_fd_sc_hd__o22a_1 _6913_ (.A1(net184),
    .A2(_0601_),
    .B1(_0602_),
    .B2(net185),
    .X(_3271_));
 sky130_fd_sc_hd__a2bb2o_1 _6914_ (.A1_N(\ann.ReLU_out[6][22] ),
    .A2_N(_0578_),
    .B1(net185),
    .B2(_0602_),
    .X(_3272_));
 sky130_fd_sc_hd__nand2_1 _6915_ (.A(_0578_),
    .B(\ann.ReLU_out[6][22] ),
    .Y(_3273_));
 sky130_fd_sc_hd__nor2_1 _6916_ (.A(_0579_),
    .B(\ann.ReLU_out[6][21] ),
    .Y(_3274_));
 sky130_fd_sc_hd__a22o_1 _6917_ (.A1(_0579_),
    .A2(\ann.ReLU_out[6][21] ),
    .B1(\ann.ReLU_out[6][20] ),
    .B2(_0580_),
    .X(_3275_));
 sky130_fd_sc_hd__nand2b_1 _6918_ (.A_N(_3274_),
    .B(_3275_),
    .Y(_3276_));
 sky130_fd_sc_hd__a21o_1 _6919_ (.A1(_3273_),
    .A2(_3276_),
    .B1(_3272_),
    .X(_3277_));
 sky130_fd_sc_hd__a21o_1 _6920_ (.A1(_3271_),
    .A2(_3277_),
    .B1(_3270_),
    .X(_3278_));
 sky130_fd_sc_hd__a21oi_1 _6921_ (.A1(_3269_),
    .A2(_3278_),
    .B1(_3268_),
    .Y(_3279_));
 sky130_fd_sc_hd__o22a_1 _6922_ (.A1(_0569_),
    .A2(\ann.ReLU_out[6][29] ),
    .B1(\ann.ReLU_out[6][28] ),
    .B2(_0571_),
    .X(_3280_));
 sky130_fd_sc_hd__and2_1 _6923_ (.A(_0569_),
    .B(\ann.ReLU_out[6][29] ),
    .X(_3281_));
 sky130_fd_sc_hd__a21oi_1 _6924_ (.A1(_0571_),
    .A2(\ann.ReLU_out[6][28] ),
    .B1(_3281_),
    .Y(_3282_));
 sky130_fd_sc_hd__o211ai_1 _6925_ (.A1(\ann.temp[27] ),
    .A2(_0598_),
    .B1(_3280_),
    .C1(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__o22a_1 _6926_ (.A1(_3280_),
    .A2(_3281_),
    .B1(_3283_),
    .B2(_3279_),
    .X(_3284_));
 sky130_fd_sc_hd__o22a_1 _6927_ (.A1(net103),
    .A2(\ann.ReLU_out[6][15] ),
    .B1(\ann.ReLU_out[6][14] ),
    .B2(net102),
    .X(_3285_));
 sky130_fd_sc_hd__a22o_1 _6928_ (.A1(net102),
    .A2(\ann.ReLU_out[6][14] ),
    .B1(\ann.ReLU_out[6][13] ),
    .B2(net101),
    .X(_3286_));
 sky130_fd_sc_hd__o22a_1 _6929_ (.A1(net101),
    .A2(\ann.ReLU_out[6][13] ),
    .B1(\ann.ReLU_out[6][12] ),
    .B2(net100),
    .X(_3287_));
 sky130_fd_sc_hd__a22o_1 _6930_ (.A1(\ann.temp[11] ),
    .A2(_0682_),
    .B1(_0683_),
    .B2(\ann.temp[10] ),
    .X(_3288_));
 sky130_fd_sc_hd__a22o_1 _6931_ (.A1(\ann.temp[9] ),
    .A2(_0684_),
    .B1(_0685_),
    .B2(net189),
    .X(_3289_));
 sky130_fd_sc_hd__o22a_1 _6932_ (.A1(\ann.temp[10] ),
    .A2(_0683_),
    .B1(_0684_),
    .B2(\ann.temp[9] ),
    .X(_3290_));
 sky130_fd_sc_hd__a21o_1 _6933_ (.A1(_3289_),
    .A2(_3290_),
    .B1(_3288_),
    .X(_3291_));
 sky130_fd_sc_hd__o2bb2a_1 _6934_ (.A1_N(net100),
    .A2_N(\ann.ReLU_out[6][12] ),
    .B1(_0682_),
    .B2(\ann.temp[11] ),
    .X(_3292_));
 sky130_fd_sc_hd__nand2_1 _6935_ (.A(_3291_),
    .B(_3292_),
    .Y(_3293_));
 sky130_fd_sc_hd__a21o_1 _6936_ (.A1(_3287_),
    .A2(_3293_),
    .B1(_3286_),
    .X(_3294_));
 sky130_fd_sc_hd__a22o_1 _6937_ (.A1(net103),
    .A2(\ann.ReLU_out[6][15] ),
    .B1(_3285_),
    .B2(_3294_),
    .X(_3295_));
 sky130_fd_sc_hd__or2_1 _6938_ (.A(net98),
    .B(\ann.ReLU_out[6][6] ),
    .X(_3296_));
 sky130_fd_sc_hd__or2_1 _6939_ (.A(net93),
    .B(\ann.ReLU_out[6][1] ),
    .X(_3297_));
 sky130_fd_sc_hd__a22o_1 _6940_ (.A1(net94),
    .A2(\ann.ReLU_out[6][2] ),
    .B1(\ann.ReLU_out[6][1] ),
    .B2(net93),
    .X(_3298_));
 sky130_fd_sc_hd__a31o_1 _6941_ (.A1(_0661_),
    .A2(\ann.ReLU_out[6][0] ),
    .A3(_3297_),
    .B1(_3298_),
    .X(_3299_));
 sky130_fd_sc_hd__o221a_1 _6942_ (.A1(net95),
    .A2(\ann.ReLU_out[6][3] ),
    .B1(\ann.ReLU_out[6][2] ),
    .B2(net94),
    .C1(_3299_),
    .X(_3300_));
 sky130_fd_sc_hd__a221o_1 _6943_ (.A1(net96),
    .A2(\ann.ReLU_out[6][4] ),
    .B1(\ann.ReLU_out[6][3] ),
    .B2(net95),
    .C1(_3300_),
    .X(_3301_));
 sky130_fd_sc_hd__o221a_1 _6944_ (.A1(net97),
    .A2(\ann.ReLU_out[6][5] ),
    .B1(\ann.ReLU_out[6][4] ),
    .B2(net96),
    .C1(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__a221o_1 _6945_ (.A1(net98),
    .A2(\ann.ReLU_out[6][6] ),
    .B1(\ann.ReLU_out[6][5] ),
    .B2(net97),
    .C1(_3302_),
    .X(_3303_));
 sky130_fd_sc_hd__a22o_1 _6946_ (.A1(net99),
    .A2(\ann.ReLU_out[6][7] ),
    .B1(_3296_),
    .B2(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__o21a_1 _6947_ (.A1(net99),
    .A2(\ann.ReLU_out[6][7] ),
    .B1(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__or4bb_1 _6948_ (.A(_3288_),
    .B(_3289_),
    .C_N(_3290_),
    .D_N(_3292_),
    .X(_3306_));
 sky130_fd_sc_hd__o221a_1 _6949_ (.A1(\ann.temp[15] ),
    .A2(_0681_),
    .B1(_0685_),
    .B2(net189),
    .C1(_3285_),
    .X(_3307_));
 sky130_fd_sc_hd__nand3b_1 _6950_ (.A_N(_3286_),
    .B(_3287_),
    .C(_3307_),
    .Y(_3308_));
 sky130_fd_sc_hd__o31a_1 _6951_ (.A1(_3305_),
    .A2(_3306_),
    .A3(_3308_),
    .B1(_3295_),
    .X(_3309_));
 sky130_fd_sc_hd__o22a_1 _6952_ (.A1(net187),
    .A2(_0678_),
    .B1(_0679_),
    .B2(net188),
    .X(_3310_));
 sky130_fd_sc_hd__nand2_1 _6953_ (.A(net187),
    .B(_0678_),
    .Y(_3311_));
 sky130_fd_sc_hd__o211ai_1 _6954_ (.A1(\ann.temp[16] ),
    .A2(_0680_),
    .B1(_3310_),
    .C1(_3311_),
    .Y(_3312_));
 sky130_fd_sc_hd__a22o_1 _6955_ (.A1(net188),
    .A2(_0679_),
    .B1(_0680_),
    .B2(\ann.temp[16] ),
    .X(_3313_));
 sky130_fd_sc_hd__xor2_1 _6956_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[6][19] ),
    .X(_3314_));
 sky130_fd_sc_hd__or4_1 _6957_ (.A(_3309_),
    .B(_3312_),
    .C(_3313_),
    .D(_3314_),
    .X(_3315_));
 sky130_fd_sc_hd__nand2_1 _6958_ (.A(_3310_),
    .B(_3313_),
    .Y(_3316_));
 sky130_fd_sc_hd__a21o_1 _6959_ (.A1(_3311_),
    .A2(_3316_),
    .B1(_3314_),
    .X(_3317_));
 sky130_fd_sc_hd__or4b_1 _6960_ (.A(_3267_),
    .B(_3268_),
    .C(_3270_),
    .D_N(_3273_),
    .X(_3318_));
 sky130_fd_sc_hd__a221o_1 _6961_ (.A1(\ann.temp[20] ),
    .A2(_0603_),
    .B1(\ann.temp[19] ),
    .B2(_0677_),
    .C1(_3283_),
    .X(_3319_));
 sky130_fd_sc_hd__or4b_1 _6962_ (.A(_3274_),
    .B(_3318_),
    .C(_3319_),
    .D_N(_3269_),
    .X(_3320_));
 sky130_fd_sc_hd__nor3_1 _6963_ (.A(_3272_),
    .B(_3275_),
    .C(_3320_),
    .Y(_3321_));
 sky130_fd_sc_hd__a41o_1 _6964_ (.A1(_3271_),
    .A2(_3315_),
    .A3(_3317_),
    .A4(_3321_),
    .B1(_3284_),
    .X(_3322_));
 sky130_fd_sc_hd__nand2_1 _6965_ (.A(\ann.temp[30] ),
    .B(_0597_),
    .Y(_3323_));
 sky130_fd_sc_hd__a21o_1 _6966_ (.A1(_3322_),
    .A2(_3323_),
    .B1(_3267_),
    .X(_3324_));
 sky130_fd_sc_hd__o22a_1 _6967_ (.A1(net103),
    .A2(\ann.ReLU_out[5][15] ),
    .B1(\ann.ReLU_out[5][14] ),
    .B2(net102),
    .X(_3325_));
 sky130_fd_sc_hd__a22o_1 _6968_ (.A1(net102),
    .A2(\ann.ReLU_out[5][14] ),
    .B1(\ann.ReLU_out[5][13] ),
    .B2(net101),
    .X(_3326_));
 sky130_fd_sc_hd__o22ai_1 _6969_ (.A1(net101),
    .A2(\ann.ReLU_out[5][13] ),
    .B1(\ann.ReLU_out[5][12] ),
    .B2(_0649_),
    .Y(_3327_));
 sky130_fd_sc_hd__o22ai_1 _6970_ (.A1(_0650_),
    .A2(\ann.ReLU_out[5][11] ),
    .B1(\ann.ReLU_out[5][10] ),
    .B2(_0651_),
    .Y(_3328_));
 sky130_fd_sc_hd__a2bb2o_1 _6971_ (.A1_N(_0652_),
    .A2_N(\ann.ReLU_out[5][9] ),
    .B1(_0676_),
    .B2(net189),
    .X(_3329_));
 sky130_fd_sc_hd__a22o_1 _6972_ (.A1(_0651_),
    .A2(\ann.ReLU_out[5][10] ),
    .B1(\ann.ReLU_out[5][9] ),
    .B2(_0652_),
    .X(_3330_));
 sky130_fd_sc_hd__and2b_1 _6973_ (.A_N(_3330_),
    .B(_3329_),
    .X(_3331_));
 sky130_fd_sc_hd__a22o_1 _6974_ (.A1(_0649_),
    .A2(\ann.ReLU_out[5][12] ),
    .B1(\ann.ReLU_out[5][11] ),
    .B2(_0650_),
    .X(_3332_));
 sky130_fd_sc_hd__o21ba_1 _6975_ (.A1(_3328_),
    .A2(_3331_),
    .B1_N(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__o21bai_1 _6976_ (.A1(_3327_),
    .A2(_3333_),
    .B1_N(_3326_),
    .Y(_3334_));
 sky130_fd_sc_hd__a22o_1 _6977_ (.A1(net103),
    .A2(\ann.ReLU_out[5][15] ),
    .B1(_3325_),
    .B2(_3334_),
    .X(_3335_));
 sky130_fd_sc_hd__or2_1 _6978_ (.A(_0655_),
    .B(\ann.ReLU_out[5][6] ),
    .X(_3336_));
 sky130_fd_sc_hd__or2_1 _6979_ (.A(net93),
    .B(\ann.ReLU_out[5][1] ),
    .X(_3337_));
 sky130_fd_sc_hd__a22o_1 _6980_ (.A1(net94),
    .A2(\ann.ReLU_out[5][2] ),
    .B1(\ann.ReLU_out[5][1] ),
    .B2(_0660_),
    .X(_3338_));
 sky130_fd_sc_hd__a31o_1 _6981_ (.A1(_0661_),
    .A2(\ann.ReLU_out[5][0] ),
    .A3(_3337_),
    .B1(_3338_),
    .X(_3339_));
 sky130_fd_sc_hd__o221a_1 _6982_ (.A1(net95),
    .A2(\ann.ReLU_out[5][3] ),
    .B1(\ann.ReLU_out[5][2] ),
    .B2(net94),
    .C1(_3339_),
    .X(_3340_));
 sky130_fd_sc_hd__a221o_1 _6983_ (.A1(net96),
    .A2(\ann.ReLU_out[5][4] ),
    .B1(\ann.ReLU_out[5][3] ),
    .B2(net95),
    .C1(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__o221a_1 _6984_ (.A1(net97),
    .A2(\ann.ReLU_out[5][5] ),
    .B1(\ann.ReLU_out[5][4] ),
    .B2(_0657_),
    .C1(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__a221o_1 _6985_ (.A1(_0655_),
    .A2(\ann.ReLU_out[5][6] ),
    .B1(\ann.ReLU_out[5][5] ),
    .B2(_0656_),
    .C1(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__a22o_1 _6986_ (.A1(net99),
    .A2(\ann.ReLU_out[5][7] ),
    .B1(_3336_),
    .B2(_3343_),
    .X(_3344_));
 sky130_fd_sc_hd__o21a_1 _6987_ (.A1(_0654_),
    .A2(\ann.ReLU_out[5][7] ),
    .B1(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__or4_1 _6988_ (.A(_3328_),
    .B(_3329_),
    .C(_3330_),
    .D(_3332_),
    .X(_3346_));
 sky130_fd_sc_hd__o221a_1 _6989_ (.A1(\ann.temp[15] ),
    .A2(_0675_),
    .B1(_0676_),
    .B2(net189),
    .C1(_3325_),
    .X(_3347_));
 sky130_fd_sc_hd__or4b_1 _6990_ (.A(_3326_),
    .B(_3327_),
    .C(_3346_),
    .D_N(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__o21a_1 _6991_ (.A1(_3345_),
    .A2(_3348_),
    .B1(_3335_),
    .X(_3349_));
 sky130_fd_sc_hd__xor2_1 _6992_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[5][19] ),
    .X(_3350_));
 sky130_fd_sc_hd__a221o_1 _6993_ (.A1(net187),
    .A2(_0673_),
    .B1(\ann.ReLU_out[5][16] ),
    .B2(_0643_),
    .C1(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__a2bb2o_1 _6994_ (.A1_N(\ann.ReLU_out[5][16] ),
    .A2_N(_0643_),
    .B1(net188),
    .B2(_0674_),
    .X(_3352_));
 sky130_fd_sc_hd__o22a_1 _6995_ (.A1(net187),
    .A2(_0673_),
    .B1(_0674_),
    .B2(net188),
    .X(_3353_));
 sky130_fd_sc_hd__or4b_1 _6996_ (.A(_3349_),
    .B(_3351_),
    .C(_3352_),
    .D_N(_3353_),
    .X(_3354_));
 sky130_fd_sc_hd__o2bb2a_1 _6997_ (.A1_N(_3352_),
    .A2_N(_3353_),
    .B1(_0640_),
    .B2(\ann.ReLU_out[5][18] ),
    .X(_3355_));
 sky130_fd_sc_hd__or2_1 _6998_ (.A(_3350_),
    .B(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__a22o_1 _6999_ (.A1(net183),
    .A2(_0608_),
    .B1(_0609_),
    .B2(net184),
    .X(_3357_));
 sky130_fd_sc_hd__o22a_1 _7000_ (.A1(net184),
    .A2(_0609_),
    .B1(_0610_),
    .B2(net185),
    .X(_3358_));
 sky130_fd_sc_hd__nand2b_1 _7001_ (.A_N(_3357_),
    .B(_3358_),
    .Y(_3359_));
 sky130_fd_sc_hd__a22o_1 _7002_ (.A1(net185),
    .A2(_0610_),
    .B1(_0611_),
    .B2(net186),
    .X(_3360_));
 sky130_fd_sc_hd__a22o_1 _7003_ (.A1(_0579_),
    .A2(\ann.ReLU_out[5][21] ),
    .B1(\ann.ReLU_out[5][20] ),
    .B2(_0580_),
    .X(_3361_));
 sky130_fd_sc_hd__a22o_1 _7004_ (.A1(\ann.temp[29] ),
    .A2(_0604_),
    .B1(_0605_),
    .B2(\ann.temp[28] ),
    .X(_3362_));
 sky130_fd_sc_hd__nor2_1 _7005_ (.A(net104),
    .B(\ann.ReLU_out[5][30] ),
    .Y(_3363_));
 sky130_fd_sc_hd__nand2_1 _7006_ (.A(net104),
    .B(\ann.ReLU_out[5][30] ),
    .Y(_3364_));
 sky130_fd_sc_hd__a22o_1 _7007_ (.A1(\ann.temp[27] ),
    .A2(_0606_),
    .B1(_0607_),
    .B2(net182),
    .X(_3365_));
 sky130_fd_sc_hd__nor2_1 _7008_ (.A(\ann.temp[29] ),
    .B(_0604_),
    .Y(_3366_));
 sky130_fd_sc_hd__nor2_1 _7009_ (.A(net186),
    .B(_0611_),
    .Y(_3367_));
 sky130_fd_sc_hd__nor2_1 _7010_ (.A(net182),
    .B(_0607_),
    .Y(_3368_));
 sky130_fd_sc_hd__or2_1 _7011_ (.A(_0579_),
    .B(\ann.ReLU_out[5][21] ),
    .X(_3369_));
 sky130_fd_sc_hd__or4b_1 _7012_ (.A(_3363_),
    .B(_3367_),
    .C(_3368_),
    .D_N(_3369_),
    .X(_3370_));
 sky130_fd_sc_hd__a221o_1 _7013_ (.A1(_0572_),
    .A2(\ann.ReLU_out[5][27] ),
    .B1(\ann.ReLU_out[5][25] ),
    .B2(_0574_),
    .C1(_3365_),
    .X(_3371_));
 sky130_fd_sc_hd__a211o_1 _7014_ (.A1(_0571_),
    .A2(\ann.ReLU_out[5][28] ),
    .B1(_3362_),
    .C1(_3366_),
    .X(_3372_));
 sky130_fd_sc_hd__o221a_1 _7015_ (.A1(_0580_),
    .A2(\ann.ReLU_out[5][20] ),
    .B1(_0639_),
    .B2(\ann.ReLU_out[5][19] ),
    .C1(_3364_),
    .X(_3373_));
 sky130_fd_sc_hd__or4b_1 _7016_ (.A(_3370_),
    .B(_3371_),
    .C(_3372_),
    .D_N(_3373_),
    .X(_3374_));
 sky130_fd_sc_hd__nor4_1 _7017_ (.A(_3359_),
    .B(_3360_),
    .C(_3361_),
    .D(_3374_),
    .Y(_3375_));
 sky130_fd_sc_hd__a21oi_1 _7018_ (.A1(_3361_),
    .A2(_3369_),
    .B1(_3367_),
    .Y(_3376_));
 sky130_fd_sc_hd__o21a_1 _7019_ (.A1(_3360_),
    .A2(_3376_),
    .B1(_3358_),
    .X(_3377_));
 sky130_fd_sc_hd__or2_1 _7020_ (.A(_3357_),
    .B(_3377_),
    .X(_3378_));
 sky130_fd_sc_hd__o221a_1 _7021_ (.A1(net182),
    .A2(_0607_),
    .B1(_0608_),
    .B2(net183),
    .C1(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__or2_1 _7022_ (.A(_3365_),
    .B(_3379_),
    .X(_3380_));
 sky130_fd_sc_hd__o221a_1 _7023_ (.A1(\ann.temp[28] ),
    .A2(_0605_),
    .B1(_0606_),
    .B2(\ann.temp[27] ),
    .C1(_3380_),
    .X(_3381_));
 sky130_fd_sc_hd__o21ba_1 _7024_ (.A1(_3362_),
    .A2(_3381_),
    .B1_N(_3366_),
    .X(_3382_));
 sky130_fd_sc_hd__o21ai_1 _7025_ (.A1(_3363_),
    .A2(_3382_),
    .B1(_3364_),
    .Y(_3383_));
 sky130_fd_sc_hd__a31o_2 _7026_ (.A1(_3354_),
    .A2(_3356_),
    .A3(_3375_),
    .B1(_3383_),
    .X(_3384_));
 sky130_fd_sc_hd__o22a_1 _7027_ (.A1(net103),
    .A2(\ann.ReLU_out[4][15] ),
    .B1(net616),
    .B2(net102),
    .X(_3385_));
 sky130_fd_sc_hd__a22o_1 _7028_ (.A1(net102),
    .A2(net616),
    .B1(\ann.ReLU_out[4][13] ),
    .B2(net101),
    .X(_3386_));
 sky130_fd_sc_hd__o22ai_1 _7029_ (.A1(net101),
    .A2(\ann.ReLU_out[4][13] ),
    .B1(\ann.ReLU_out[4][12] ),
    .B2(net100),
    .Y(_3387_));
 sky130_fd_sc_hd__o22ai_1 _7030_ (.A1(_0650_),
    .A2(\ann.ReLU_out[4][11] ),
    .B1(\ann.ReLU_out[4][10] ),
    .B2(_0651_),
    .Y(_3388_));
 sky130_fd_sc_hd__a2bb2o_1 _7031_ (.A1_N(_0652_),
    .A2_N(\ann.ReLU_out[4][9] ),
    .B1(_0672_),
    .B2(net189),
    .X(_3389_));
 sky130_fd_sc_hd__a22o_1 _7032_ (.A1(_0651_),
    .A2(\ann.ReLU_out[4][10] ),
    .B1(\ann.ReLU_out[4][9] ),
    .B2(_0652_),
    .X(_3390_));
 sky130_fd_sc_hd__and2b_1 _7033_ (.A_N(_3390_),
    .B(_3389_),
    .X(_3391_));
 sky130_fd_sc_hd__a22o_1 _7034_ (.A1(net100),
    .A2(\ann.ReLU_out[4][12] ),
    .B1(\ann.ReLU_out[4][11] ),
    .B2(_0650_),
    .X(_3392_));
 sky130_fd_sc_hd__o21ba_1 _7035_ (.A1(_3388_),
    .A2(_3391_),
    .B1_N(_3392_),
    .X(_3393_));
 sky130_fd_sc_hd__o21bai_1 _7036_ (.A1(_3387_),
    .A2(_3393_),
    .B1_N(_3386_),
    .Y(_3394_));
 sky130_fd_sc_hd__a22o_1 _7037_ (.A1(net103),
    .A2(\ann.ReLU_out[4][15] ),
    .B1(_3385_),
    .B2(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__or2_1 _7038_ (.A(net98),
    .B(\ann.ReLU_out[4][6] ),
    .X(_3396_));
 sky130_fd_sc_hd__or2_1 _7039_ (.A(_0660_),
    .B(\ann.ReLU_out[4][1] ),
    .X(_3397_));
 sky130_fd_sc_hd__a22o_1 _7040_ (.A1(net94),
    .A2(\ann.ReLU_out[4][2] ),
    .B1(\ann.ReLU_out[4][1] ),
    .B2(net93),
    .X(_3398_));
 sky130_fd_sc_hd__a31o_1 _7041_ (.A1(_0661_),
    .A2(\ann.ReLU_out[4][0] ),
    .A3(_3397_),
    .B1(_3398_),
    .X(_3399_));
 sky130_fd_sc_hd__o221a_1 _7042_ (.A1(net95),
    .A2(\ann.ReLU_out[4][3] ),
    .B1(\ann.ReLU_out[4][2] ),
    .B2(_0659_),
    .C1(_3399_),
    .X(_3400_));
 sky130_fd_sc_hd__a221o_1 _7043_ (.A1(net96),
    .A2(\ann.ReLU_out[4][4] ),
    .B1(\ann.ReLU_out[4][3] ),
    .B2(_0658_),
    .C1(_3400_),
    .X(_3401_));
 sky130_fd_sc_hd__o221a_1 _7044_ (.A1(net97),
    .A2(\ann.ReLU_out[4][5] ),
    .B1(\ann.ReLU_out[4][4] ),
    .B2(_0657_),
    .C1(_3401_),
    .X(_3402_));
 sky130_fd_sc_hd__a221o_1 _7045_ (.A1(net98),
    .A2(\ann.ReLU_out[4][6] ),
    .B1(\ann.ReLU_out[4][5] ),
    .B2(net97),
    .C1(_3402_),
    .X(_3403_));
 sky130_fd_sc_hd__a22o_1 _7046_ (.A1(net99),
    .A2(\ann.ReLU_out[4][7] ),
    .B1(_3396_),
    .B2(_3403_),
    .X(_3404_));
 sky130_fd_sc_hd__o21a_1 _7047_ (.A1(_0654_),
    .A2(\ann.ReLU_out[4][7] ),
    .B1(_3404_),
    .X(_3405_));
 sky130_fd_sc_hd__or4_1 _7048_ (.A(_3388_),
    .B(_3389_),
    .C(_3390_),
    .D(_3392_),
    .X(_3406_));
 sky130_fd_sc_hd__o221a_1 _7049_ (.A1(\ann.temp[15] ),
    .A2(_0671_),
    .B1(_0672_),
    .B2(net189),
    .C1(_3385_),
    .X(_3407_));
 sky130_fd_sc_hd__or4b_1 _7050_ (.A(_3386_),
    .B(_3387_),
    .C(_3406_),
    .D_N(_3407_),
    .X(_3408_));
 sky130_fd_sc_hd__o21a_1 _7051_ (.A1(_3405_),
    .A2(_3408_),
    .B1(_3395_),
    .X(_3409_));
 sky130_fd_sc_hd__xor2_1 _7052_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[4][19] ),
    .X(_3410_));
 sky130_fd_sc_hd__a221o_1 _7053_ (.A1(net187),
    .A2(_0669_),
    .B1(\ann.ReLU_out[4][16] ),
    .B2(_0643_),
    .C1(_3410_),
    .X(_3411_));
 sky130_fd_sc_hd__a2bb2o_1 _7054_ (.A1_N(\ann.ReLU_out[4][16] ),
    .A2_N(_0643_),
    .B1(net188),
    .B2(_0670_),
    .X(_3412_));
 sky130_fd_sc_hd__o22a_1 _7055_ (.A1(net187),
    .A2(_0669_),
    .B1(_0670_),
    .B2(net188),
    .X(_3413_));
 sky130_fd_sc_hd__or4b_1 _7056_ (.A(_3409_),
    .B(_3411_),
    .C(_3412_),
    .D_N(_3413_),
    .X(_3414_));
 sky130_fd_sc_hd__o2bb2a_1 _7057_ (.A1_N(_3412_),
    .A2_N(_3413_),
    .B1(_0640_),
    .B2(net603),
    .X(_3415_));
 sky130_fd_sc_hd__or2_1 _7058_ (.A(_3410_),
    .B(_3415_),
    .X(_3416_));
 sky130_fd_sc_hd__a22o_1 _7059_ (.A1(net183),
    .A2(_0616_),
    .B1(_0617_),
    .B2(net184),
    .X(_3417_));
 sky130_fd_sc_hd__o22a_1 _7060_ (.A1(net184),
    .A2(_0617_),
    .B1(_0618_),
    .B2(\ann.temp[23] ),
    .X(_3418_));
 sky130_fd_sc_hd__nand2b_1 _7061_ (.A_N(_3417_),
    .B(_3418_),
    .Y(_3419_));
 sky130_fd_sc_hd__a22o_1 _7062_ (.A1(\ann.temp[23] ),
    .A2(_0618_),
    .B1(_0619_),
    .B2(net186),
    .X(_3420_));
 sky130_fd_sc_hd__a22o_1 _7063_ (.A1(_0579_),
    .A2(\ann.ReLU_out[4][21] ),
    .B1(net589),
    .B2(_0580_),
    .X(_3421_));
 sky130_fd_sc_hd__a22o_1 _7064_ (.A1(\ann.temp[29] ),
    .A2(_0612_),
    .B1(_0613_),
    .B2(\ann.temp[28] ),
    .X(_3422_));
 sky130_fd_sc_hd__nor2_1 _7065_ (.A(net104),
    .B(\ann.ReLU_out[4][30] ),
    .Y(_3423_));
 sky130_fd_sc_hd__nand2_1 _7066_ (.A(net104),
    .B(\ann.ReLU_out[4][30] ),
    .Y(_3424_));
 sky130_fd_sc_hd__a22o_1 _7067_ (.A1(\ann.temp[27] ),
    .A2(_0614_),
    .B1(_0615_),
    .B2(net182),
    .X(_3425_));
 sky130_fd_sc_hd__nor2_1 _7068_ (.A(\ann.temp[29] ),
    .B(_0612_),
    .Y(_3426_));
 sky130_fd_sc_hd__nor2_1 _7069_ (.A(net186),
    .B(_0619_),
    .Y(_3427_));
 sky130_fd_sc_hd__nor2_1 _7070_ (.A(net182),
    .B(_0615_),
    .Y(_3428_));
 sky130_fd_sc_hd__or2_1 _7071_ (.A(_0579_),
    .B(\ann.ReLU_out[4][21] ),
    .X(_3429_));
 sky130_fd_sc_hd__or4b_1 _7072_ (.A(_3423_),
    .B(_3427_),
    .C(_3428_),
    .D_N(_3429_),
    .X(_3430_));
 sky130_fd_sc_hd__a221o_1 _7073_ (.A1(_0572_),
    .A2(\ann.ReLU_out[4][27] ),
    .B1(\ann.ReLU_out[4][25] ),
    .B2(_0574_),
    .C1(_3425_),
    .X(_3431_));
 sky130_fd_sc_hd__a211o_1 _7074_ (.A1(_0571_),
    .A2(net674),
    .B1(_3422_),
    .C1(_3426_),
    .X(_3432_));
 sky130_fd_sc_hd__o221a_1 _7075_ (.A1(_0580_),
    .A2(\ann.ReLU_out[4][20] ),
    .B1(_0639_),
    .B2(\ann.ReLU_out[4][19] ),
    .C1(_3424_),
    .X(_3433_));
 sky130_fd_sc_hd__or4b_1 _7076_ (.A(_3430_),
    .B(_3431_),
    .C(_3432_),
    .D_N(_3433_),
    .X(_3434_));
 sky130_fd_sc_hd__nor4_2 _7077_ (.A(_3419_),
    .B(_3420_),
    .C(_3421_),
    .D(_3434_),
    .Y(_3435_));
 sky130_fd_sc_hd__a21oi_1 _7078_ (.A1(_3421_),
    .A2(_3429_),
    .B1(_3427_),
    .Y(_3436_));
 sky130_fd_sc_hd__o21a_1 _7079_ (.A1(_3420_),
    .A2(_3436_),
    .B1(_3418_),
    .X(_3437_));
 sky130_fd_sc_hd__or2_1 _7080_ (.A(_3417_),
    .B(_3437_),
    .X(_3438_));
 sky130_fd_sc_hd__o221a_1 _7081_ (.A1(net182),
    .A2(_0615_),
    .B1(_0616_),
    .B2(net183),
    .C1(_3438_),
    .X(_3439_));
 sky130_fd_sc_hd__or2_1 _7082_ (.A(_3425_),
    .B(_3439_),
    .X(_3440_));
 sky130_fd_sc_hd__o221a_1 _7083_ (.A1(\ann.temp[28] ),
    .A2(_0613_),
    .B1(_0614_),
    .B2(\ann.temp[27] ),
    .C1(_3440_),
    .X(_3441_));
 sky130_fd_sc_hd__o21ba_1 _7084_ (.A1(_3422_),
    .A2(_3441_),
    .B1_N(_3426_),
    .X(_3442_));
 sky130_fd_sc_hd__o21ai_1 _7085_ (.A1(_3423_),
    .A2(_3442_),
    .B1(_3424_),
    .Y(_3443_));
 sky130_fd_sc_hd__a31o_2 _7086_ (.A1(_3414_),
    .A2(_3416_),
    .A3(_3435_),
    .B1(_3443_),
    .X(_3444_));
 sky130_fd_sc_hd__and2_1 _7087_ (.A(net104),
    .B(\ann.ReLU_out[3][30] ),
    .X(_3445_));
 sky130_fd_sc_hd__o2bb2a_1 _7088_ (.A1_N(_0573_),
    .A2_N(\ann.ReLU_out[3][26] ),
    .B1(_0620_),
    .B2(net183),
    .X(_3446_));
 sky130_fd_sc_hd__a22o_1 _7089_ (.A1(net183),
    .A2(_0620_),
    .B1(_0621_),
    .B2(net184),
    .X(_3447_));
 sky130_fd_sc_hd__o22a_1 _7090_ (.A1(net184),
    .A2(_0621_),
    .B1(_0622_),
    .B2(\ann.temp[23] ),
    .X(_3448_));
 sky130_fd_sc_hd__inv_2 _7091_ (.A(_3448_),
    .Y(_3449_));
 sky130_fd_sc_hd__a22o_1 _7092_ (.A1(net185),
    .A2(_0622_),
    .B1(_0623_),
    .B2(\ann.temp[22] ),
    .X(_3450_));
 sky130_fd_sc_hd__nor2_1 _7093_ (.A(net186),
    .B(_0623_),
    .Y(_3451_));
 sky130_fd_sc_hd__a22o_1 _7094_ (.A1(_0579_),
    .A2(\ann.ReLU_out[3][21] ),
    .B1(\ann.ReLU_out[3][20] ),
    .B2(_0580_),
    .X(_3452_));
 sky130_fd_sc_hd__or2_1 _7095_ (.A(_0579_),
    .B(\ann.ReLU_out[3][21] ),
    .X(_3453_));
 sky130_fd_sc_hd__a21oi_1 _7096_ (.A1(_3452_),
    .A2(_3453_),
    .B1(_3451_),
    .Y(_3454_));
 sky130_fd_sc_hd__o21a_1 _7097_ (.A1(_3450_),
    .A2(_3454_),
    .B1(_3448_),
    .X(_3455_));
 sky130_fd_sc_hd__o21ai_1 _7098_ (.A1(_3447_),
    .A2(_3455_),
    .B1(_3446_),
    .Y(_3456_));
 sky130_fd_sc_hd__o221a_1 _7099_ (.A1(_0572_),
    .A2(\ann.ReLU_out[3][27] ),
    .B1(\ann.ReLU_out[3][26] ),
    .B2(_0573_),
    .C1(_3456_),
    .X(_3457_));
 sky130_fd_sc_hd__or2_1 _7100_ (.A(_0569_),
    .B(\ann.ReLU_out[3][29] ),
    .X(_3458_));
 sky130_fd_sc_hd__o21ai_1 _7101_ (.A1(_0571_),
    .A2(net645),
    .B1(_3458_),
    .Y(_3459_));
 sky130_fd_sc_hd__and2_1 _7102_ (.A(_0569_),
    .B(\ann.ReLU_out[3][29] ),
    .X(_3460_));
 sky130_fd_sc_hd__a211o_1 _7103_ (.A1(_0571_),
    .A2(net645),
    .B1(_3459_),
    .C1(_3460_),
    .X(_3461_));
 sky130_fd_sc_hd__and2_1 _7104_ (.A(_0572_),
    .B(\ann.ReLU_out[3][27] ),
    .X(_3462_));
 sky130_fd_sc_hd__or2_1 _7105_ (.A(net104),
    .B(\ann.ReLU_out[3][30] ),
    .X(_3463_));
 sky130_fd_sc_hd__o311a_1 _7106_ (.A1(_0571_),
    .A2(net645),
    .A3(_3460_),
    .B1(_3463_),
    .C1(_3458_),
    .X(_3464_));
 sky130_fd_sc_hd__o31a_1 _7107_ (.A1(_3457_),
    .A2(_3461_),
    .A3(_3462_),
    .B1(_3464_),
    .X(_3465_));
 sky130_fd_sc_hd__o22a_1 _7108_ (.A1(net103),
    .A2(\ann.ReLU_out[3][15] ),
    .B1(\ann.ReLU_out[3][14] ),
    .B2(net102),
    .X(_3466_));
 sky130_fd_sc_hd__a22o_1 _7109_ (.A1(net102),
    .A2(\ann.ReLU_out[3][14] ),
    .B1(\ann.ReLU_out[3][13] ),
    .B2(net101),
    .X(_3467_));
 sky130_fd_sc_hd__o22ai_1 _7110_ (.A1(net101),
    .A2(\ann.ReLU_out[3][13] ),
    .B1(\ann.ReLU_out[3][12] ),
    .B2(net100),
    .Y(_3468_));
 sky130_fd_sc_hd__o22ai_1 _7111_ (.A1(_0650_),
    .A2(\ann.ReLU_out[3][11] ),
    .B1(\ann.ReLU_out[3][10] ),
    .B2(_0651_),
    .Y(_3469_));
 sky130_fd_sc_hd__a2bb2o_1 _7112_ (.A1_N(_0652_),
    .A2_N(\ann.ReLU_out[3][9] ),
    .B1(_0668_),
    .B2(net189),
    .X(_3470_));
 sky130_fd_sc_hd__a22o_1 _7113_ (.A1(_0651_),
    .A2(\ann.ReLU_out[3][10] ),
    .B1(\ann.ReLU_out[3][9] ),
    .B2(_0652_),
    .X(_3471_));
 sky130_fd_sc_hd__and2b_1 _7114_ (.A_N(_3471_),
    .B(_3470_),
    .X(_3472_));
 sky130_fd_sc_hd__a22o_1 _7115_ (.A1(net100),
    .A2(\ann.ReLU_out[3][12] ),
    .B1(\ann.ReLU_out[3][11] ),
    .B2(_0650_),
    .X(_3473_));
 sky130_fd_sc_hd__o21ba_1 _7116_ (.A1(_3469_),
    .A2(_3472_),
    .B1_N(_3473_),
    .X(_3474_));
 sky130_fd_sc_hd__nor2_1 _7117_ (.A(_3468_),
    .B(_3474_),
    .Y(_3475_));
 sky130_fd_sc_hd__o21a_1 _7118_ (.A1(_3467_),
    .A2(_3475_),
    .B1(_3466_),
    .X(_3476_));
 sky130_fd_sc_hd__a21oi_1 _7119_ (.A1(net103),
    .A2(\ann.ReLU_out[3][15] ),
    .B1(_3476_),
    .Y(_3477_));
 sky130_fd_sc_hd__or2_1 _7120_ (.A(net98),
    .B(\ann.ReLU_out[3][6] ),
    .X(_3478_));
 sky130_fd_sc_hd__or2_1 _7121_ (.A(net93),
    .B(\ann.ReLU_out[3][1] ),
    .X(_3479_));
 sky130_fd_sc_hd__a22o_1 _7122_ (.A1(net94),
    .A2(\ann.ReLU_out[3][2] ),
    .B1(\ann.ReLU_out[3][1] ),
    .B2(net93),
    .X(_3480_));
 sky130_fd_sc_hd__a31o_1 _7123_ (.A1(_0661_),
    .A2(\ann.ReLU_out[3][0] ),
    .A3(_3479_),
    .B1(_3480_),
    .X(_3481_));
 sky130_fd_sc_hd__o221a_1 _7124_ (.A1(net95),
    .A2(\ann.ReLU_out[3][3] ),
    .B1(\ann.ReLU_out[3][2] ),
    .B2(net94),
    .C1(_3481_),
    .X(_3482_));
 sky130_fd_sc_hd__a221o_1 _7125_ (.A1(net96),
    .A2(\ann.ReLU_out[3][4] ),
    .B1(\ann.ReLU_out[3][3] ),
    .B2(net95),
    .C1(_3482_),
    .X(_3483_));
 sky130_fd_sc_hd__o221a_1 _7126_ (.A1(net97),
    .A2(\ann.ReLU_out[3][5] ),
    .B1(\ann.ReLU_out[3][4] ),
    .B2(net96),
    .C1(_3483_),
    .X(_3484_));
 sky130_fd_sc_hd__a221o_1 _7127_ (.A1(net98),
    .A2(\ann.ReLU_out[3][6] ),
    .B1(\ann.ReLU_out[3][5] ),
    .B2(net97),
    .C1(_3484_),
    .X(_3485_));
 sky130_fd_sc_hd__a22o_1 _7128_ (.A1(net99),
    .A2(\ann.ReLU_out[3][7] ),
    .B1(_3478_),
    .B2(_3485_),
    .X(_3486_));
 sky130_fd_sc_hd__o21a_1 _7129_ (.A1(net99),
    .A2(\ann.ReLU_out[3][7] ),
    .B1(_3486_),
    .X(_3487_));
 sky130_fd_sc_hd__or4_1 _7130_ (.A(_3469_),
    .B(_3470_),
    .C(_3471_),
    .D(_3473_),
    .X(_3488_));
 sky130_fd_sc_hd__o221a_1 _7131_ (.A1(\ann.temp[15] ),
    .A2(_0667_),
    .B1(_0668_),
    .B2(net189),
    .C1(_3466_),
    .X(_3489_));
 sky130_fd_sc_hd__or4b_1 _7132_ (.A(_3467_),
    .B(_3468_),
    .C(_3488_),
    .D_N(_3489_),
    .X(_3490_));
 sky130_fd_sc_hd__nor2_1 _7133_ (.A(_3487_),
    .B(_3490_),
    .Y(_3491_));
 sky130_fd_sc_hd__o22a_1 _7134_ (.A1(_0642_),
    .A2(\ann.ReLU_out[3][17] ),
    .B1(\ann.ReLU_out[3][16] ),
    .B2(_0643_),
    .X(_3492_));
 sky130_fd_sc_hd__nand2_1 _7135_ (.A(net187),
    .B(_0666_),
    .Y(_3493_));
 sky130_fd_sc_hd__o2bb2a_1 _7136_ (.A1_N(\ann.ReLU_out[3][17] ),
    .A2_N(_0642_),
    .B1(net187),
    .B2(_0666_),
    .X(_3494_));
 sky130_fd_sc_hd__xor2_1 _7137_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[3][19] ),
    .X(_3495_));
 sky130_fd_sc_hd__a221oi_1 _7138_ (.A1(net187),
    .A2(_0666_),
    .B1(\ann.ReLU_out[3][16] ),
    .B2(_0643_),
    .C1(_3495_),
    .Y(_3496_));
 sky130_fd_sc_hd__o2111a_1 _7139_ (.A1(_3477_),
    .A2(_3491_),
    .B1(_3492_),
    .C1(_3494_),
    .D1(_3496_),
    .X(_3497_));
 sky130_fd_sc_hd__or4_1 _7140_ (.A(_3447_),
    .B(_3449_),
    .C(_3450_),
    .D(_3452_),
    .X(_3498_));
 sky130_fd_sc_hd__o221ai_1 _7141_ (.A1(_0572_),
    .A2(\ann.ReLU_out[3][27] ),
    .B1(\ann.ReLU_out[3][26] ),
    .B2(_0573_),
    .C1(_3446_),
    .Y(_3499_));
 sky130_fd_sc_hd__or4b_1 _7142_ (.A(_3445_),
    .B(_3451_),
    .C(_3462_),
    .D_N(_3463_),
    .X(_3500_));
 sky130_fd_sc_hd__o221a_1 _7143_ (.A1(_0580_),
    .A2(\ann.ReLU_out[3][20] ),
    .B1(_0639_),
    .B2(\ann.ReLU_out[3][19] ),
    .C1(_3453_),
    .X(_3501_));
 sky130_fd_sc_hd__or4b_1 _7144_ (.A(_3498_),
    .B(_3499_),
    .C(_3500_),
    .D_N(_3501_),
    .X(_3502_));
 sky130_fd_sc_hd__nand2b_1 _7145_ (.A_N(_3492_),
    .B(_3494_),
    .Y(_3503_));
 sky130_fd_sc_hd__a21oi_1 _7146_ (.A1(_3493_),
    .A2(_3503_),
    .B1(_3495_),
    .Y(_3504_));
 sky130_fd_sc_hd__or4_1 _7147_ (.A(_3461_),
    .B(_3497_),
    .C(_3502_),
    .D(_3504_),
    .X(_3505_));
 sky130_fd_sc_hd__or3b_1 _7148_ (.A(_3445_),
    .B(_3465_),
    .C_N(_3505_),
    .X(_3506_));
 sky130_fd_sc_hd__inv_2 _7149_ (.A(_3506_),
    .Y(_3507_));
 sky130_fd_sc_hd__o22a_1 _7150_ (.A1(net103),
    .A2(\ann.ReLU_out[2][15] ),
    .B1(\ann.ReLU_out[2][14] ),
    .B2(net102),
    .X(_3508_));
 sky130_fd_sc_hd__a22o_1 _7151_ (.A1(net102),
    .A2(\ann.ReLU_out[2][14] ),
    .B1(\ann.ReLU_out[2][13] ),
    .B2(net101),
    .X(_3509_));
 sky130_fd_sc_hd__o22ai_1 _7152_ (.A1(_0648_),
    .A2(\ann.ReLU_out[2][13] ),
    .B1(\ann.ReLU_out[2][12] ),
    .B2(net100),
    .Y(_3510_));
 sky130_fd_sc_hd__o22ai_1 _7153_ (.A1(_0650_),
    .A2(\ann.ReLU_out[2][11] ),
    .B1(\ann.ReLU_out[2][10] ),
    .B2(_0651_),
    .Y(_3511_));
 sky130_fd_sc_hd__a2bb2o_1 _7154_ (.A1_N(_0652_),
    .A2_N(\ann.ReLU_out[2][9] ),
    .B1(_0665_),
    .B2(net189),
    .X(_3512_));
 sky130_fd_sc_hd__a22o_1 _7155_ (.A1(_0651_),
    .A2(\ann.ReLU_out[2][10] ),
    .B1(\ann.ReLU_out[2][9] ),
    .B2(_0652_),
    .X(_3513_));
 sky130_fd_sc_hd__and2b_1 _7156_ (.A_N(_3513_),
    .B(_3512_),
    .X(_3514_));
 sky130_fd_sc_hd__a22o_1 _7157_ (.A1(net100),
    .A2(\ann.ReLU_out[2][12] ),
    .B1(\ann.ReLU_out[2][11] ),
    .B2(_0650_),
    .X(_3515_));
 sky130_fd_sc_hd__o21ba_1 _7158_ (.A1(_3511_),
    .A2(_3514_),
    .B1_N(_3515_),
    .X(_3516_));
 sky130_fd_sc_hd__o21bai_1 _7159_ (.A1(_3510_),
    .A2(_3516_),
    .B1_N(_3509_),
    .Y(_3517_));
 sky130_fd_sc_hd__a22o_1 _7160_ (.A1(net103),
    .A2(net695),
    .B1(_3508_),
    .B2(_3517_),
    .X(_3518_));
 sky130_fd_sc_hd__or2_1 _7161_ (.A(net98),
    .B(\ann.ReLU_out[2][6] ),
    .X(_3519_));
 sky130_fd_sc_hd__or2_1 _7162_ (.A(net93),
    .B(\ann.ReLU_out[2][1] ),
    .X(_3520_));
 sky130_fd_sc_hd__a22o_1 _7163_ (.A1(net94),
    .A2(\ann.ReLU_out[2][2] ),
    .B1(\ann.ReLU_out[2][1] ),
    .B2(net93),
    .X(_3521_));
 sky130_fd_sc_hd__a31o_1 _7164_ (.A1(_0661_),
    .A2(\ann.ReLU_out[2][0] ),
    .A3(_3520_),
    .B1(_3521_),
    .X(_3522_));
 sky130_fd_sc_hd__o221a_1 _7165_ (.A1(net95),
    .A2(\ann.ReLU_out[2][3] ),
    .B1(\ann.ReLU_out[2][2] ),
    .B2(net94),
    .C1(_3522_),
    .X(_3523_));
 sky130_fd_sc_hd__a221o_1 _7166_ (.A1(net96),
    .A2(\ann.ReLU_out[2][4] ),
    .B1(\ann.ReLU_out[2][3] ),
    .B2(_0658_),
    .C1(_3523_),
    .X(_3524_));
 sky130_fd_sc_hd__o221a_1 _7167_ (.A1(net97),
    .A2(\ann.ReLU_out[2][5] ),
    .B1(\ann.ReLU_out[2][4] ),
    .B2(net96),
    .C1(_3524_),
    .X(_3525_));
 sky130_fd_sc_hd__a221o_1 _7168_ (.A1(net98),
    .A2(\ann.ReLU_out[2][6] ),
    .B1(\ann.ReLU_out[2][5] ),
    .B2(net97),
    .C1(_3525_),
    .X(_3526_));
 sky130_fd_sc_hd__a22o_1 _7169_ (.A1(net99),
    .A2(\ann.ReLU_out[2][7] ),
    .B1(_3519_),
    .B2(_3526_),
    .X(_3527_));
 sky130_fd_sc_hd__o21a_1 _7170_ (.A1(net99),
    .A2(\ann.ReLU_out[2][7] ),
    .B1(_3527_),
    .X(_3528_));
 sky130_fd_sc_hd__or4_1 _7171_ (.A(_3511_),
    .B(_3512_),
    .C(_3513_),
    .D(_3515_),
    .X(_3529_));
 sky130_fd_sc_hd__o221a_1 _7172_ (.A1(\ann.temp[15] ),
    .A2(_0664_),
    .B1(_0665_),
    .B2(\ann.temp[8] ),
    .C1(_3508_),
    .X(_3530_));
 sky130_fd_sc_hd__or4b_1 _7173_ (.A(_3509_),
    .B(_3510_),
    .C(_3529_),
    .D_N(_3530_),
    .X(_3531_));
 sky130_fd_sc_hd__o21a_1 _7174_ (.A1(_3528_),
    .A2(_3531_),
    .B1(_3518_),
    .X(_3532_));
 sky130_fd_sc_hd__xor2_1 _7175_ (.A(\ann.temp[19] ),
    .B(\ann.ReLU_out[2][19] ),
    .X(_3533_));
 sky130_fd_sc_hd__a221o_1 _7176_ (.A1(net187),
    .A2(_0662_),
    .B1(\ann.ReLU_out[2][16] ),
    .B2(_0643_),
    .C1(_3533_),
    .X(_3534_));
 sky130_fd_sc_hd__a2bb2o_1 _7177_ (.A1_N(\ann.ReLU_out[2][16] ),
    .A2_N(_0643_),
    .B1(net188),
    .B2(_0663_),
    .X(_3535_));
 sky130_fd_sc_hd__o22a_1 _7178_ (.A1(\ann.temp[18] ),
    .A2(_0662_),
    .B1(_0663_),
    .B2(net188),
    .X(_3536_));
 sky130_fd_sc_hd__or4b_1 _7179_ (.A(_3532_),
    .B(_3534_),
    .C(_3535_),
    .D_N(_3536_),
    .X(_3537_));
 sky130_fd_sc_hd__o2bb2a_1 _7180_ (.A1_N(_3535_),
    .A2_N(_3536_),
    .B1(_0640_),
    .B2(\ann.ReLU_out[2][18] ),
    .X(_3538_));
 sky130_fd_sc_hd__a22o_1 _7181_ (.A1(net183),
    .A2(_0628_),
    .B1(_0629_),
    .B2(net184),
    .X(_3539_));
 sky130_fd_sc_hd__o22a_1 _7182_ (.A1(\ann.temp[24] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(net185),
    .X(_3540_));
 sky130_fd_sc_hd__nand2b_1 _7183_ (.A_N(_3539_),
    .B(_3540_),
    .Y(_3541_));
 sky130_fd_sc_hd__a22o_1 _7184_ (.A1(net185),
    .A2(_0630_),
    .B1(_0631_),
    .B2(\ann.temp[22] ),
    .X(_3542_));
 sky130_fd_sc_hd__a22o_1 _7185_ (.A1(_0579_),
    .A2(net639),
    .B1(\ann.ReLU_out[2][20] ),
    .B2(_0580_),
    .X(_3543_));
 sky130_fd_sc_hd__a22o_1 _7186_ (.A1(\ann.temp[29] ),
    .A2(_0624_),
    .B1(_0625_),
    .B2(\ann.temp[28] ),
    .X(_3544_));
 sky130_fd_sc_hd__nor2_1 _7187_ (.A(net104),
    .B(\ann.ReLU_out[2][30] ),
    .Y(_3545_));
 sky130_fd_sc_hd__nand2_1 _7188_ (.A(net104),
    .B(\ann.ReLU_out[2][30] ),
    .Y(_3546_));
 sky130_fd_sc_hd__a22o_1 _7189_ (.A1(\ann.temp[27] ),
    .A2(_0626_),
    .B1(_0627_),
    .B2(net182),
    .X(_3547_));
 sky130_fd_sc_hd__nor2_1 _7190_ (.A(\ann.temp[29] ),
    .B(_0624_),
    .Y(_3548_));
 sky130_fd_sc_hd__nor2_1 _7191_ (.A(\ann.temp[22] ),
    .B(_0631_),
    .Y(_3549_));
 sky130_fd_sc_hd__nor2_1 _7192_ (.A(net182),
    .B(_0627_),
    .Y(_3550_));
 sky130_fd_sc_hd__or2_1 _7193_ (.A(_0579_),
    .B(\ann.ReLU_out[2][21] ),
    .X(_3551_));
 sky130_fd_sc_hd__or4b_1 _7194_ (.A(_3545_),
    .B(_3549_),
    .C(_3550_),
    .D_N(_3551_),
    .X(_3552_));
 sky130_fd_sc_hd__a221o_1 _7195_ (.A1(_0572_),
    .A2(\ann.ReLU_out[2][27] ),
    .B1(\ann.ReLU_out[2][25] ),
    .B2(_0574_),
    .C1(_3547_),
    .X(_3553_));
 sky130_fd_sc_hd__a211o_1 _7196_ (.A1(_0571_),
    .A2(net618),
    .B1(_3544_),
    .C1(_3548_),
    .X(_3554_));
 sky130_fd_sc_hd__o221a_1 _7197_ (.A1(_0580_),
    .A2(\ann.ReLU_out[2][20] ),
    .B1(_0639_),
    .B2(\ann.ReLU_out[2][19] ),
    .C1(_3546_),
    .X(_3555_));
 sky130_fd_sc_hd__or4b_1 _7198_ (.A(_3552_),
    .B(_3553_),
    .C(_3554_),
    .D_N(_3555_),
    .X(_3556_));
 sky130_fd_sc_hd__nor4_1 _7199_ (.A(_3541_),
    .B(_3542_),
    .C(_3543_),
    .D(_3556_),
    .Y(_3557_));
 sky130_fd_sc_hd__o211ai_1 _7200_ (.A1(_3533_),
    .A2(_3538_),
    .B1(_3557_),
    .C1(_3537_),
    .Y(_3558_));
 sky130_fd_sc_hd__a21oi_1 _7201_ (.A1(_3543_),
    .A2(_3551_),
    .B1(_3549_),
    .Y(_3559_));
 sky130_fd_sc_hd__o21a_1 _7202_ (.A1(_3542_),
    .A2(_3559_),
    .B1(_3540_),
    .X(_3560_));
 sky130_fd_sc_hd__or2_1 _7203_ (.A(_3539_),
    .B(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__o221a_1 _7204_ (.A1(\ann.temp[26] ),
    .A2(_0627_),
    .B1(_0628_),
    .B2(net183),
    .C1(_3561_),
    .X(_3562_));
 sky130_fd_sc_hd__or2_1 _7205_ (.A(_3547_),
    .B(_3562_),
    .X(_3563_));
 sky130_fd_sc_hd__o221a_1 _7206_ (.A1(\ann.temp[28] ),
    .A2(_0625_),
    .B1(_0626_),
    .B2(\ann.temp[27] ),
    .C1(_3563_),
    .X(_3564_));
 sky130_fd_sc_hd__o21ba_1 _7207_ (.A1(_3544_),
    .A2(_3564_),
    .B1_N(_3548_),
    .X(_3565_));
 sky130_fd_sc_hd__o211a_2 _7208_ (.A1(_3545_),
    .A2(_3565_),
    .B1(_3558_),
    .C1(_3546_),
    .X(_3566_));
 sky130_fd_sc_hd__o22a_1 _7209_ (.A1(\ann.ReLU_out[1][15] ),
    .A2(_0646_),
    .B1(\ann.ReLU_out[1][14] ),
    .B2(_0647_),
    .X(_3567_));
 sky130_fd_sc_hd__a22o_1 _7210_ (.A1(\ann.ReLU_out[1][14] ),
    .A2(_0647_),
    .B1(\ann.ReLU_out[1][13] ),
    .B2(_0648_),
    .X(_3568_));
 sky130_fd_sc_hd__o22ai_2 _7211_ (.A1(\ann.ReLU_out[1][13] ),
    .A2(_0648_),
    .B1(net100),
    .B2(\ann.ReLU_out[1][12] ),
    .Y(_3569_));
 sky130_fd_sc_hd__o22ai_1 _7212_ (.A1(\ann.ReLU_out[1][11] ),
    .A2(_0650_),
    .B1(\ann.ReLU_out[1][10] ),
    .B2(_0651_),
    .Y(_3570_));
 sky130_fd_sc_hd__a2bb2o_1 _7213_ (.A1_N(\ann.ReLU_out[1][9] ),
    .A2_N(_0652_),
    .B1(\ann.temp[8] ),
    .B2(_0653_),
    .X(_3571_));
 sky130_fd_sc_hd__a22o_1 _7214_ (.A1(\ann.ReLU_out[1][10] ),
    .A2(_0651_),
    .B1(\ann.ReLU_out[1][9] ),
    .B2(_0652_),
    .X(_3572_));
 sky130_fd_sc_hd__and2b_1 _7215_ (.A_N(_3572_),
    .B(_3571_),
    .X(_3573_));
 sky130_fd_sc_hd__a22o_1 _7216_ (.A1(_0649_),
    .A2(\ann.ReLU_out[1][12] ),
    .B1(\ann.ReLU_out[1][11] ),
    .B2(_0650_),
    .X(_3574_));
 sky130_fd_sc_hd__o21ba_1 _7217_ (.A1(_3570_),
    .A2(_3573_),
    .B1_N(_3574_),
    .X(_3575_));
 sky130_fd_sc_hd__o21bai_1 _7218_ (.A1(_3569_),
    .A2(_3575_),
    .B1_N(_3568_),
    .Y(_3576_));
 sky130_fd_sc_hd__a22o_1 _7219_ (.A1(\ann.ReLU_out[1][15] ),
    .A2(_0646_),
    .B1(_3567_),
    .B2(_3576_),
    .X(_3577_));
 sky130_fd_sc_hd__or2_1 _7220_ (.A(\ann.ReLU_out[1][6] ),
    .B(net98),
    .X(_3578_));
 sky130_fd_sc_hd__or2_1 _7221_ (.A(\ann.ReLU_out[1][1] ),
    .B(net93),
    .X(_3579_));
 sky130_fd_sc_hd__a22o_1 _7222_ (.A1(\ann.ReLU_out[1][2] ),
    .A2(_0659_),
    .B1(\ann.ReLU_out[1][1] ),
    .B2(net93),
    .X(_3580_));
 sky130_fd_sc_hd__a31o_1 _7223_ (.A1(\ann.ReLU_out[1][0] ),
    .A2(_0661_),
    .A3(_3579_),
    .B1(_3580_),
    .X(_3581_));
 sky130_fd_sc_hd__o221a_1 _7224_ (.A1(\ann.ReLU_out[1][3] ),
    .A2(net95),
    .B1(\ann.ReLU_out[1][2] ),
    .B2(net94),
    .C1(_3581_),
    .X(_3582_));
 sky130_fd_sc_hd__a221o_1 _7225_ (.A1(net96),
    .A2(\ann.ReLU_out[1][4] ),
    .B1(\ann.ReLU_out[1][3] ),
    .B2(net95),
    .C1(_3582_),
    .X(_3583_));
 sky130_fd_sc_hd__o221a_1 _7226_ (.A1(\ann.ReLU_out[1][5] ),
    .A2(net97),
    .B1(net96),
    .B2(\ann.ReLU_out[1][4] ),
    .C1(_3583_),
    .X(_3584_));
 sky130_fd_sc_hd__a221o_1 _7227_ (.A1(\ann.ReLU_out[1][6] ),
    .A2(net98),
    .B1(\ann.ReLU_out[1][5] ),
    .B2(_0656_),
    .C1(_3584_),
    .X(_3585_));
 sky130_fd_sc_hd__a22o_1 _7228_ (.A1(\ann.ReLU_out[1][7] ),
    .A2(net99),
    .B1(_3578_),
    .B2(_3585_),
    .X(_3586_));
 sky130_fd_sc_hd__o21a_1 _7229_ (.A1(\ann.ReLU_out[1][7] ),
    .A2(net99),
    .B1(_3586_),
    .X(_3587_));
 sky130_fd_sc_hd__or4_1 _7230_ (.A(_3570_),
    .B(_3571_),
    .C(_3572_),
    .D(_3574_),
    .X(_3588_));
 sky130_fd_sc_hd__o221a_1 _7231_ (.A1(_0645_),
    .A2(\ann.temp[15] ),
    .B1(\ann.temp[8] ),
    .B2(_0653_),
    .C1(_3567_),
    .X(_3589_));
 sky130_fd_sc_hd__or4b_1 _7232_ (.A(_3568_),
    .B(_3569_),
    .C(_3588_),
    .D_N(_3589_),
    .X(_3590_));
 sky130_fd_sc_hd__o21a_1 _7233_ (.A1(_3587_),
    .A2(_3590_),
    .B1(_3577_),
    .X(_3591_));
 sky130_fd_sc_hd__a22o_1 _7234_ (.A1(_0641_),
    .A2(\ann.temp[17] ),
    .B1(\ann.temp[16] ),
    .B2(_0644_),
    .X(_3592_));
 sky130_fd_sc_hd__or2_1 _7235_ (.A(\ann.ReLU_out[1][18] ),
    .B(_0640_),
    .X(_3593_));
 sky130_fd_sc_hd__o21ai_1 _7236_ (.A1(\ann.temp[16] ),
    .A2(_0644_),
    .B1(_3593_),
    .Y(_3594_));
 sky130_fd_sc_hd__o2bb2a_1 _7237_ (.A1_N(\ann.ReLU_out[1][18] ),
    .A2_N(_0640_),
    .B1(_0641_),
    .B2(\ann.temp[17] ),
    .X(_3595_));
 sky130_fd_sc_hd__or2_1 _7238_ (.A(\ann.ReLU_out[1][19] ),
    .B(_0639_),
    .X(_3596_));
 sky130_fd_sc_hd__nand2_1 _7239_ (.A(\ann.ReLU_out[1][19] ),
    .B(_0639_),
    .Y(_3597_));
 sky130_fd_sc_hd__nand2_1 _7240_ (.A(_3596_),
    .B(_3597_),
    .Y(_3598_));
 sky130_fd_sc_hd__and2b_1 _7241_ (.A_N(_3592_),
    .B(_3595_),
    .X(_3599_));
 sky130_fd_sc_hd__or4b_1 _7242_ (.A(_3591_),
    .B(_3594_),
    .C(_3598_),
    .D_N(_3599_),
    .X(_3600_));
 sky130_fd_sc_hd__a22o_1 _7243_ (.A1(\ann.temp[23] ),
    .A2(_0637_),
    .B1(_0638_),
    .B2(net186),
    .X(_3601_));
 sky130_fd_sc_hd__a22o_1 _7244_ (.A1(_0579_),
    .A2(net648),
    .B1(\ann.ReLU_out[1][20] ),
    .B2(_0580_),
    .X(_3602_));
 sky130_fd_sc_hd__a22o_1 _7245_ (.A1(net183),
    .A2(_0635_),
    .B1(_0636_),
    .B2(\ann.temp[24] ),
    .X(_3603_));
 sky130_fd_sc_hd__o22a_1 _7246_ (.A1(net184),
    .A2(_0636_),
    .B1(_0637_),
    .B2(\ann.temp[23] ),
    .X(_3604_));
 sky130_fd_sc_hd__nor4b_1 _7247_ (.A(_3601_),
    .B(_3602_),
    .C(_3603_),
    .D_N(_3604_),
    .Y(_3605_));
 sky130_fd_sc_hd__a22o_1 _7248_ (.A1(\ann.temp[27] ),
    .A2(_0633_),
    .B1(_0634_),
    .B2(\ann.temp[26] ),
    .X(_3606_));
 sky130_fd_sc_hd__o22a_1 _7249_ (.A1(\ann.temp[26] ),
    .A2(_0634_),
    .B1(_0635_),
    .B2(net183),
    .X(_3607_));
 sky130_fd_sc_hd__or2_1 _7250_ (.A(_0579_),
    .B(\ann.ReLU_out[1][21] ),
    .X(_3608_));
 sky130_fd_sc_hd__nor2_1 _7251_ (.A(net104),
    .B(\ann.ReLU_out[1][30] ),
    .Y(_3609_));
 sky130_fd_sc_hd__nor2_1 _7252_ (.A(_0571_),
    .B(\ann.ReLU_out[1][28] ),
    .Y(_3610_));
 sky130_fd_sc_hd__nor2_1 _7253_ (.A(_0569_),
    .B(\ann.ReLU_out[1][29] ),
    .Y(_3611_));
 sky130_fd_sc_hd__nand2_1 _7254_ (.A(_0569_),
    .B(\ann.ReLU_out[1][29] ),
    .Y(_3612_));
 sky130_fd_sc_hd__a22o_1 _7255_ (.A1(_0569_),
    .A2(\ann.ReLU_out[1][29] ),
    .B1(\ann.ReLU_out[1][28] ),
    .B2(_0571_),
    .X(_3613_));
 sky130_fd_sc_hd__nor3_1 _7256_ (.A(_3610_),
    .B(_3611_),
    .C(_3613_),
    .Y(_3614_));
 sky130_fd_sc_hd__a22o_1 _7257_ (.A1(_0567_),
    .A2(\ann.ReLU_out[1][30] ),
    .B1(\ann.ReLU_out[1][22] ),
    .B2(_0578_),
    .X(_3615_));
 sky130_fd_sc_hd__a211o_1 _7258_ (.A1(_0572_),
    .A2(\ann.ReLU_out[1][27] ),
    .B1(_3609_),
    .C1(_3615_),
    .X(_3616_));
 sky130_fd_sc_hd__nor2_1 _7259_ (.A(_3606_),
    .B(_3616_),
    .Y(_3617_));
 sky130_fd_sc_hd__o211a_1 _7260_ (.A1(_0580_),
    .A2(\ann.ReLU_out[1][20] ),
    .B1(_3596_),
    .C1(_3608_),
    .X(_3618_));
 sky130_fd_sc_hd__and4_1 _7261_ (.A(_3607_),
    .B(_3614_),
    .C(_3617_),
    .D(_3618_),
    .X(_3619_));
 sky130_fd_sc_hd__nand2_1 _7262_ (.A(_3605_),
    .B(_3619_),
    .Y(_3620_));
 sky130_fd_sc_hd__a21boi_1 _7263_ (.A1(_3592_),
    .A2(_3595_),
    .B1_N(_3593_),
    .Y(_3621_));
 sky130_fd_sc_hd__o2bb2a_1 _7264_ (.A1_N(_3602_),
    .A2_N(_3608_),
    .B1(\ann.temp[22] ),
    .B2(_0638_),
    .X(_3622_));
 sky130_fd_sc_hd__o21a_1 _7265_ (.A1(_3601_),
    .A2(_3622_),
    .B1(_3604_),
    .X(_3623_));
 sky130_fd_sc_hd__o21a_1 _7266_ (.A1(_3603_),
    .A2(_3623_),
    .B1(_3607_),
    .X(_3624_));
 sky130_fd_sc_hd__o22a_1 _7267_ (.A1(\ann.temp[27] ),
    .A2(_0633_),
    .B1(_3606_),
    .B2(_3624_),
    .X(_3625_));
 sky130_fd_sc_hd__or2_1 _7268_ (.A(_3609_),
    .B(_3611_),
    .X(_3626_));
 sky130_fd_sc_hd__a221o_1 _7269_ (.A1(_3610_),
    .A2(_3612_),
    .B1(_3614_),
    .B2(_3625_),
    .C1(_3626_),
    .X(_3627_));
 sky130_fd_sc_hd__o21ai_1 _7270_ (.A1(_3598_),
    .A2(_3621_),
    .B1(_3600_),
    .Y(_3628_));
 sky130_fd_sc_hd__o221a_2 _7271_ (.A1(\ann.temp[30] ),
    .A2(_0632_),
    .B1(_3620_),
    .B2(_3628_),
    .C1(_3627_),
    .X(_3629_));
 sky130_fd_sc_hd__inv_2 _7272_ (.A(net41),
    .Y(_3630_));
 sky130_fd_sc_hd__a21oi_1 _7273_ (.A1(net43),
    .A2(_3630_),
    .B1(_3506_),
    .Y(_3631_));
 sky130_fd_sc_hd__o21ba_1 _7274_ (.A1(net54),
    .A2(_3631_),
    .B1_N(net56),
    .X(_3632_));
 sky130_fd_sc_hd__o21bai_1 _7275_ (.A1(net44),
    .A2(_3632_),
    .B1_N(net48),
    .Y(_3633_));
 sky130_fd_sc_hd__a21bo_1 _7276_ (.A1(net50),
    .A2(_3633_),
    .B1_N(net38),
    .X(_0100_));
 sky130_fd_sc_hd__and2_2 _7277_ (.A(net38),
    .B(net50),
    .X(_3634_));
 sky130_fd_sc_hd__clkinv_4 _7278_ (.A(_3634_),
    .Y(_0103_));
 sky130_fd_sc_hd__or2_2 _7279_ (.A(net56),
    .B(net53),
    .X(_3635_));
 sky130_fd_sc_hd__a21oi_2 _7280_ (.A1(net36),
    .A2(net42),
    .B1(_3635_),
    .Y(_3636_));
 sky130_fd_sc_hd__o31a_4 _7281_ (.A1(net48),
    .A2(net44),
    .A3(_3636_),
    .B1(_3634_),
    .X(_0101_));
 sky130_fd_sc_hd__o31a_4 _7282_ (.A1(net47),
    .A2(net44),
    .A3(_3635_),
    .B1(_3634_),
    .X(_0102_));
 sky130_fd_sc_hd__and2_2 _7283_ (.A(net210),
    .B(net19),
    .X(_3637_));
 sky130_fd_sc_hd__mux2_1 _7284_ (.A0(\ann.ReLU_out[1][0] ),
    .A1(\ann.ReLU_out[0][0] ),
    .S(net41),
    .X(_3638_));
 sky130_fd_sc_hd__mux2_1 _7285_ (.A0(\ann.ReLU_out[2][0] ),
    .A1(_3638_),
    .S(net43),
    .X(_3639_));
 sky130_fd_sc_hd__mux2_1 _7286_ (.A0(\ann.ReLU_out[3][0] ),
    .A1(_3639_),
    .S(net37),
    .X(_3640_));
 sky130_fd_sc_hd__mux2_1 _7287_ (.A0(_3640_),
    .A1(\ann.ReLU_out[4][0] ),
    .S(net54),
    .X(_3641_));
 sky130_fd_sc_hd__mux2_1 _7288_ (.A0(_3641_),
    .A1(net347),
    .S(net56),
    .X(_3642_));
 sky130_fd_sc_hd__mux2_1 _7289_ (.A0(_3642_),
    .A1(\ann.ReLU_out[6][0] ),
    .S(net46),
    .X(_3643_));
 sky130_fd_sc_hd__mux2_1 _7290_ (.A0(_3643_),
    .A1(\ann.ReLU_out[7][0] ),
    .S(net49),
    .X(_3644_));
 sky130_fd_sc_hd__mux2_1 _7291_ (.A0(\ann.ReLU_out[8][0] ),
    .A1(_3644_),
    .S(net52),
    .X(_3645_));
 sky130_fd_sc_hd__mux2_1 _7292_ (.A0(\ann.ReLU_out[9][0] ),
    .A1(_3645_),
    .S(_3142_),
    .X(_3646_));
 sky130_fd_sc_hd__mux2_1 _7293_ (.A0(net353),
    .A1(_3646_),
    .S(net90),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _7294_ (.A0(\ann.ReLU_out[1][1] ),
    .A1(\ann.ReLU_out[0][1] ),
    .S(net41),
    .X(_3647_));
 sky130_fd_sc_hd__mux2_1 _7295_ (.A0(\ann.ReLU_out[2][1] ),
    .A1(_3647_),
    .S(net43),
    .X(_3648_));
 sky130_fd_sc_hd__mux2_1 _7296_ (.A0(\ann.ReLU_out[3][1] ),
    .A1(_3648_),
    .S(net37),
    .X(_3649_));
 sky130_fd_sc_hd__mux2_1 _7297_ (.A0(_3649_),
    .A1(\ann.ReLU_out[4][1] ),
    .S(_3444_),
    .X(_3650_));
 sky130_fd_sc_hd__mux2_1 _7298_ (.A0(_3650_),
    .A1(\ann.ReLU_out[5][1] ),
    .S(_3384_),
    .X(_3651_));
 sky130_fd_sc_hd__mux2_1 _7299_ (.A0(_3651_),
    .A1(\ann.ReLU_out[6][1] ),
    .S(net46),
    .X(_3652_));
 sky130_fd_sc_hd__mux2_1 _7300_ (.A0(_3652_),
    .A1(\ann.ReLU_out[7][1] ),
    .S(net49),
    .X(_3653_));
 sky130_fd_sc_hd__mux2_1 _7301_ (.A0(\ann.ReLU_out[8][1] ),
    .A1(_3653_),
    .S(net52),
    .X(_3654_));
 sky130_fd_sc_hd__mux2_1 _7302_ (.A0(\ann.ReLU_out[9][1] ),
    .A1(_3654_),
    .S(_3142_),
    .X(_3655_));
 sky130_fd_sc_hd__mux2_1 _7303_ (.A0(net365),
    .A1(_3655_),
    .S(net90),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _7304_ (.A0(\ann.ReLU_out[1][2] ),
    .A1(\ann.ReLU_out[0][2] ),
    .S(net41),
    .X(_3656_));
 sky130_fd_sc_hd__mux2_1 _7305_ (.A0(\ann.ReLU_out[2][2] ),
    .A1(_3656_),
    .S(net43),
    .X(_3657_));
 sky130_fd_sc_hd__mux2_1 _7306_ (.A0(\ann.ReLU_out[3][2] ),
    .A1(_3657_),
    .S(net37),
    .X(_3658_));
 sky130_fd_sc_hd__mux2_1 _7307_ (.A0(_3658_),
    .A1(\ann.ReLU_out[4][2] ),
    .S(net54),
    .X(_3659_));
 sky130_fd_sc_hd__mux2_1 _7308_ (.A0(_3659_),
    .A1(\ann.ReLU_out[5][2] ),
    .S(_3384_),
    .X(_3660_));
 sky130_fd_sc_hd__mux2_1 _7309_ (.A0(_3660_),
    .A1(\ann.ReLU_out[6][2] ),
    .S(net46),
    .X(_3661_));
 sky130_fd_sc_hd__mux2_1 _7310_ (.A0(_3661_),
    .A1(\ann.ReLU_out[7][2] ),
    .S(net49),
    .X(_3662_));
 sky130_fd_sc_hd__mux2_1 _7311_ (.A0(\ann.ReLU_out[8][2] ),
    .A1(_3662_),
    .S(net52),
    .X(_3663_));
 sky130_fd_sc_hd__mux2_1 _7312_ (.A0(\ann.ReLU_out[9][2] ),
    .A1(_3663_),
    .S(net39),
    .X(_3664_));
 sky130_fd_sc_hd__mux2_1 _7313_ (.A0(net343),
    .A1(_3664_),
    .S(net90),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _7314_ (.A0(\ann.ReLU_out[1][3] ),
    .A1(\ann.ReLU_out[0][3] ),
    .S(net41),
    .X(_3665_));
 sky130_fd_sc_hd__mux2_1 _7315_ (.A0(\ann.ReLU_out[2][3] ),
    .A1(_3665_),
    .S(net43),
    .X(_3666_));
 sky130_fd_sc_hd__mux2_1 _7316_ (.A0(\ann.ReLU_out[3][3] ),
    .A1(_3666_),
    .S(net37),
    .X(_3667_));
 sky130_fd_sc_hd__mux2_1 _7317_ (.A0(_3667_),
    .A1(\ann.ReLU_out[4][3] ),
    .S(net54),
    .X(_3668_));
 sky130_fd_sc_hd__mux2_1 _7318_ (.A0(_3668_),
    .A1(\ann.ReLU_out[5][3] ),
    .S(net56),
    .X(_3669_));
 sky130_fd_sc_hd__mux2_1 _7319_ (.A0(_3669_),
    .A1(\ann.ReLU_out[6][3] ),
    .S(net46),
    .X(_3670_));
 sky130_fd_sc_hd__mux2_1 _7320_ (.A0(_3670_),
    .A1(\ann.ReLU_out[7][3] ),
    .S(net49),
    .X(_3671_));
 sky130_fd_sc_hd__mux2_1 _7321_ (.A0(\ann.ReLU_out[8][3] ),
    .A1(_3671_),
    .S(net52),
    .X(_3672_));
 sky130_fd_sc_hd__mux2_1 _7322_ (.A0(\ann.ReLU_out[9][3] ),
    .A1(_3672_),
    .S(net39),
    .X(_3673_));
 sky130_fd_sc_hd__mux2_1 _7323_ (.A0(net349),
    .A1(_3673_),
    .S(net90),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _7324_ (.A0(\ann.ReLU_out[1][4] ),
    .A1(\ann.ReLU_out[0][4] ),
    .S(net41),
    .X(_3674_));
 sky130_fd_sc_hd__mux2_1 _7325_ (.A0(\ann.ReLU_out[2][4] ),
    .A1(_3674_),
    .S(net43),
    .X(_3675_));
 sky130_fd_sc_hd__mux2_1 _7326_ (.A0(\ann.ReLU_out[3][4] ),
    .A1(_3675_),
    .S(net37),
    .X(_3676_));
 sky130_fd_sc_hd__mux2_1 _7327_ (.A0(_3676_),
    .A1(\ann.ReLU_out[4][4] ),
    .S(net54),
    .X(_3677_));
 sky130_fd_sc_hd__mux2_1 _7328_ (.A0(_3677_),
    .A1(\ann.ReLU_out[5][4] ),
    .S(net56),
    .X(_3678_));
 sky130_fd_sc_hd__mux2_1 _7329_ (.A0(_3678_),
    .A1(\ann.ReLU_out[6][4] ),
    .S(net46),
    .X(_3679_));
 sky130_fd_sc_hd__mux2_1 _7330_ (.A0(_3679_),
    .A1(\ann.ReLU_out[7][4] ),
    .S(net49),
    .X(_3680_));
 sky130_fd_sc_hd__mux2_1 _7331_ (.A0(\ann.ReLU_out[8][4] ),
    .A1(_3680_),
    .S(net52),
    .X(_3681_));
 sky130_fd_sc_hd__mux2_1 _7332_ (.A0(\ann.ReLU_out[9][4] ),
    .A1(_3681_),
    .S(net39),
    .X(_3682_));
 sky130_fd_sc_hd__mux2_1 _7333_ (.A0(net351),
    .A1(_3682_),
    .S(net90),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _7334_ (.A0(\ann.ReLU_out[1][5] ),
    .A1(\ann.ReLU_out[0][5] ),
    .S(net41),
    .X(_3683_));
 sky130_fd_sc_hd__mux2_1 _7335_ (.A0(\ann.ReLU_out[2][5] ),
    .A1(_3683_),
    .S(net43),
    .X(_3684_));
 sky130_fd_sc_hd__mux2_1 _7336_ (.A0(\ann.ReLU_out[3][5] ),
    .A1(_3684_),
    .S(net37),
    .X(_3685_));
 sky130_fd_sc_hd__mux2_1 _7337_ (.A0(_3685_),
    .A1(\ann.ReLU_out[4][5] ),
    .S(net54),
    .X(_3686_));
 sky130_fd_sc_hd__mux2_1 _7338_ (.A0(_3686_),
    .A1(\ann.ReLU_out[5][5] ),
    .S(net56),
    .X(_3687_));
 sky130_fd_sc_hd__mux2_1 _7339_ (.A0(_3687_),
    .A1(\ann.ReLU_out[6][5] ),
    .S(net46),
    .X(_3688_));
 sky130_fd_sc_hd__mux2_1 _7340_ (.A0(_3688_),
    .A1(\ann.ReLU_out[7][5] ),
    .S(net49),
    .X(_3689_));
 sky130_fd_sc_hd__mux2_1 _7341_ (.A0(\ann.ReLU_out[8][5] ),
    .A1(_3689_),
    .S(net52),
    .X(_3690_));
 sky130_fd_sc_hd__mux2_1 _7342_ (.A0(\ann.ReLU_out[9][5] ),
    .A1(_3690_),
    .S(net39),
    .X(_3691_));
 sky130_fd_sc_hd__mux2_1 _7343_ (.A0(net329),
    .A1(_3691_),
    .S(net90),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _7344_ (.A0(\ann.ReLU_out[1][6] ),
    .A1(\ann.ReLU_out[0][6] ),
    .S(net41),
    .X(_3692_));
 sky130_fd_sc_hd__mux2_1 _7345_ (.A0(\ann.ReLU_out[2][6] ),
    .A1(_3692_),
    .S(net43),
    .X(_3693_));
 sky130_fd_sc_hd__mux2_1 _7346_ (.A0(\ann.ReLU_out[3][6] ),
    .A1(_3693_),
    .S(net37),
    .X(_3694_));
 sky130_fd_sc_hd__mux2_1 _7347_ (.A0(_3694_),
    .A1(\ann.ReLU_out[4][6] ),
    .S(net54),
    .X(_3695_));
 sky130_fd_sc_hd__mux2_1 _7348_ (.A0(_3695_),
    .A1(\ann.ReLU_out[5][6] ),
    .S(net56),
    .X(_3696_));
 sky130_fd_sc_hd__mux2_1 _7349_ (.A0(_3696_),
    .A1(\ann.ReLU_out[6][6] ),
    .S(net46),
    .X(_3697_));
 sky130_fd_sc_hd__mux2_1 _7350_ (.A0(_3697_),
    .A1(\ann.ReLU_out[7][6] ),
    .S(net49),
    .X(_3698_));
 sky130_fd_sc_hd__mux2_1 _7351_ (.A0(\ann.ReLU_out[8][6] ),
    .A1(_3698_),
    .S(net52),
    .X(_3699_));
 sky130_fd_sc_hd__mux2_1 _7352_ (.A0(\ann.ReLU_out[9][6] ),
    .A1(_3699_),
    .S(net39),
    .X(_3700_));
 sky130_fd_sc_hd__mux2_1 _7353_ (.A0(net379),
    .A1(_3700_),
    .S(net90),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _7354_ (.A0(\ann.ReLU_out[1][7] ),
    .A1(\ann.ReLU_out[0][7] ),
    .S(net41),
    .X(_3701_));
 sky130_fd_sc_hd__mux2_1 _7355_ (.A0(\ann.ReLU_out[2][7] ),
    .A1(_3701_),
    .S(_3566_),
    .X(_3702_));
 sky130_fd_sc_hd__mux2_1 _7356_ (.A0(\ann.ReLU_out[3][7] ),
    .A1(_3702_),
    .S(net37),
    .X(_3703_));
 sky130_fd_sc_hd__mux2_1 _7357_ (.A0(_3703_),
    .A1(\ann.ReLU_out[4][7] ),
    .S(net54),
    .X(_3704_));
 sky130_fd_sc_hd__mux2_1 _7358_ (.A0(_3704_),
    .A1(\ann.ReLU_out[5][7] ),
    .S(net56),
    .X(_3705_));
 sky130_fd_sc_hd__mux2_1 _7359_ (.A0(_3705_),
    .A1(\ann.ReLU_out[6][7] ),
    .S(net46),
    .X(_3706_));
 sky130_fd_sc_hd__mux2_1 _7360_ (.A0(_3706_),
    .A1(\ann.ReLU_out[7][7] ),
    .S(net49),
    .X(_3707_));
 sky130_fd_sc_hd__mux2_1 _7361_ (.A0(\ann.ReLU_out[8][7] ),
    .A1(_3707_),
    .S(net52),
    .X(_3708_));
 sky130_fd_sc_hd__mux2_1 _7362_ (.A0(\ann.ReLU_out[9][7] ),
    .A1(_3708_),
    .S(_3142_),
    .X(_3709_));
 sky130_fd_sc_hd__mux2_1 _7363_ (.A0(net333),
    .A1(_3709_),
    .S(net90),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _7364_ (.A0(\ann.ReLU_out[1][8] ),
    .A1(\ann.ReLU_out[0][8] ),
    .S(net40),
    .X(_3710_));
 sky130_fd_sc_hd__mux2_1 _7365_ (.A0(\ann.ReLU_out[2][8] ),
    .A1(_3710_),
    .S(net42),
    .X(_3711_));
 sky130_fd_sc_hd__mux2_1 _7366_ (.A0(\ann.ReLU_out[3][8] ),
    .A1(_3711_),
    .S(net36),
    .X(_3712_));
 sky130_fd_sc_hd__mux2_1 _7367_ (.A0(_3712_),
    .A1(net423),
    .S(net53),
    .X(_3713_));
 sky130_fd_sc_hd__mux2_1 _7368_ (.A0(_3713_),
    .A1(net430),
    .S(net56),
    .X(_3714_));
 sky130_fd_sc_hd__a21oi_1 _7369_ (.A1(_0685_),
    .A2(net45),
    .B1(net47),
    .Y(_3715_));
 sky130_fd_sc_hd__o21a_1 _7370_ (.A1(net45),
    .A2(_3714_),
    .B1(_3715_),
    .X(_3716_));
 sky130_fd_sc_hd__a21bo_1 _7371_ (.A1(net497),
    .A2(net48),
    .B1_N(net51),
    .X(_3717_));
 sky130_fd_sc_hd__o22a_1 _7372_ (.A1(net545),
    .A2(net50),
    .B1(_3716_),
    .B2(_3717_),
    .X(_3718_));
 sky130_fd_sc_hd__mux2_1 _7373_ (.A0(net429),
    .A1(_3718_),
    .S(net38),
    .X(_3719_));
 sky130_fd_sc_hd__mux2_1 _7374_ (.A0(net189),
    .A1(_3719_),
    .S(net89),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _7375_ (.A0(\ann.ReLU_out[1][9] ),
    .A1(\ann.ReLU_out[0][9] ),
    .S(net40),
    .X(_3720_));
 sky130_fd_sc_hd__mux2_1 _7376_ (.A0(\ann.ReLU_out[2][9] ),
    .A1(_3720_),
    .S(net42),
    .X(_3721_));
 sky130_fd_sc_hd__mux2_1 _7377_ (.A0(\ann.ReLU_out[3][9] ),
    .A1(_3721_),
    .S(net36),
    .X(_3722_));
 sky130_fd_sc_hd__mux2_1 _7378_ (.A0(_3722_),
    .A1(\ann.ReLU_out[4][9] ),
    .S(net53),
    .X(_3723_));
 sky130_fd_sc_hd__mux2_1 _7379_ (.A0(_3723_),
    .A1(net553),
    .S(net55),
    .X(_3724_));
 sky130_fd_sc_hd__mux2_1 _7380_ (.A0(_3724_),
    .A1(net488),
    .S(net45),
    .X(_3725_));
 sky130_fd_sc_hd__mux2_1 _7381_ (.A0(_3725_),
    .A1(net469),
    .S(net48),
    .X(_3726_));
 sky130_fd_sc_hd__mux2_1 _7382_ (.A0(net426),
    .A1(_3726_),
    .S(net51),
    .X(_3727_));
 sky130_fd_sc_hd__mux2_1 _7383_ (.A0(net434),
    .A1(_3727_),
    .S(net38),
    .X(_3728_));
 sky130_fd_sc_hd__mux2_1 _7384_ (.A0(net747),
    .A1(_3728_),
    .S(net89),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _7385_ (.A0(\ann.ReLU_out[1][10] ),
    .A1(\ann.ReLU_out[0][10] ),
    .S(net40),
    .X(_3729_));
 sky130_fd_sc_hd__mux2_1 _7386_ (.A0(\ann.ReLU_out[2][10] ),
    .A1(_3729_),
    .S(net42),
    .X(_3730_));
 sky130_fd_sc_hd__mux2_1 _7387_ (.A0(\ann.ReLU_out[3][10] ),
    .A1(_3730_),
    .S(net36),
    .X(_3731_));
 sky130_fd_sc_hd__mux2_1 _7388_ (.A0(_3731_),
    .A1(\ann.ReLU_out[4][10] ),
    .S(net53),
    .X(_3732_));
 sky130_fd_sc_hd__mux2_1 _7389_ (.A0(_3732_),
    .A1(\ann.ReLU_out[5][10] ),
    .S(net55),
    .X(_3733_));
 sky130_fd_sc_hd__mux2_1 _7390_ (.A0(_3733_),
    .A1(net421),
    .S(net45),
    .X(_3734_));
 sky130_fd_sc_hd__mux2_1 _7391_ (.A0(_3734_),
    .A1(net508),
    .S(net48),
    .X(_3735_));
 sky130_fd_sc_hd__mux2_1 _7392_ (.A0(net442),
    .A1(_3735_),
    .S(net51),
    .X(_3736_));
 sky130_fd_sc_hd__mux2_1 _7393_ (.A0(net510),
    .A1(_3736_),
    .S(net39),
    .X(_3737_));
 sky130_fd_sc_hd__mux2_1 _7394_ (.A0(net750),
    .A1(_3737_),
    .S(net89),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _7395_ (.A0(\ann.ReLU_out[1][11] ),
    .A1(\ann.ReLU_out[0][11] ),
    .S(net40),
    .X(_3738_));
 sky130_fd_sc_hd__mux2_1 _7396_ (.A0(\ann.ReLU_out[2][11] ),
    .A1(_3738_),
    .S(net42),
    .X(_3739_));
 sky130_fd_sc_hd__mux2_1 _7397_ (.A0(\ann.ReLU_out[3][11] ),
    .A1(_3739_),
    .S(net36),
    .X(_3740_));
 sky130_fd_sc_hd__mux2_1 _7398_ (.A0(_3740_),
    .A1(\ann.ReLU_out[4][11] ),
    .S(net53),
    .X(_3741_));
 sky130_fd_sc_hd__mux2_1 _7399_ (.A0(_3741_),
    .A1(\ann.ReLU_out[5][11] ),
    .S(net56),
    .X(_3742_));
 sky130_fd_sc_hd__mux2_1 _7400_ (.A0(_3742_),
    .A1(net484),
    .S(net45),
    .X(_3743_));
 sky130_fd_sc_hd__mux2_1 _7401_ (.A0(_3743_),
    .A1(net458),
    .S(net48),
    .X(_3744_));
 sky130_fd_sc_hd__mux2_1 _7402_ (.A0(net435),
    .A1(_3744_),
    .S(net51),
    .X(_3745_));
 sky130_fd_sc_hd__mux2_1 _7403_ (.A0(net473),
    .A1(_3745_),
    .S(net39),
    .X(_3746_));
 sky130_fd_sc_hd__mux2_1 _7404_ (.A0(net753),
    .A1(_3746_),
    .S(net89),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _7405_ (.A0(\ann.ReLU_out[1][12] ),
    .A1(\ann.ReLU_out[0][12] ),
    .S(net40),
    .X(_3747_));
 sky130_fd_sc_hd__mux2_1 _7406_ (.A0(\ann.ReLU_out[2][12] ),
    .A1(_3747_),
    .S(net42),
    .X(_3748_));
 sky130_fd_sc_hd__mux2_1 _7407_ (.A0(\ann.ReLU_out[3][12] ),
    .A1(_3748_),
    .S(net36),
    .X(_3749_));
 sky130_fd_sc_hd__mux2_1 _7408_ (.A0(_3749_),
    .A1(\ann.ReLU_out[4][12] ),
    .S(net53),
    .X(_3750_));
 sky130_fd_sc_hd__mux2_1 _7409_ (.A0(_3750_),
    .A1(\ann.ReLU_out[5][12] ),
    .S(net56),
    .X(_3751_));
 sky130_fd_sc_hd__mux2_1 _7410_ (.A0(_3751_),
    .A1(\ann.ReLU_out[6][12] ),
    .S(net45),
    .X(_3752_));
 sky130_fd_sc_hd__mux2_1 _7411_ (.A0(_3752_),
    .A1(\ann.ReLU_out[7][12] ),
    .S(net48),
    .X(_3753_));
 sky130_fd_sc_hd__mux2_1 _7412_ (.A0(\ann.ReLU_out[8][12] ),
    .A1(_3753_),
    .S(net51),
    .X(_3754_));
 sky130_fd_sc_hd__mux2_1 _7413_ (.A0(\ann.ReLU_out[9][12] ),
    .A1(_3754_),
    .S(net39),
    .X(_3755_));
 sky130_fd_sc_hd__mux2_1 _7414_ (.A0(net339),
    .A1(_3755_),
    .S(net89),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _7415_ (.A0(\ann.ReLU_out[1][13] ),
    .A1(\ann.ReLU_out[0][13] ),
    .S(net40),
    .X(_3756_));
 sky130_fd_sc_hd__mux2_1 _7416_ (.A0(\ann.ReLU_out[2][13] ),
    .A1(_3756_),
    .S(net42),
    .X(_3757_));
 sky130_fd_sc_hd__mux2_1 _7417_ (.A0(\ann.ReLU_out[3][13] ),
    .A1(_3757_),
    .S(net36),
    .X(_3758_));
 sky130_fd_sc_hd__mux2_1 _7418_ (.A0(_3758_),
    .A1(\ann.ReLU_out[4][13] ),
    .S(net54),
    .X(_3759_));
 sky130_fd_sc_hd__mux2_1 _7419_ (.A0(_3759_),
    .A1(\ann.ReLU_out[5][13] ),
    .S(net55),
    .X(_3760_));
 sky130_fd_sc_hd__mux2_1 _7420_ (.A0(_3760_),
    .A1(\ann.ReLU_out[6][13] ),
    .S(net45),
    .X(_3761_));
 sky130_fd_sc_hd__mux2_1 _7421_ (.A0(_3761_),
    .A1(\ann.ReLU_out[7][13] ),
    .S(net48),
    .X(_3762_));
 sky130_fd_sc_hd__mux2_1 _7422_ (.A0(\ann.ReLU_out[8][13] ),
    .A1(_3762_),
    .S(net51),
    .X(_3763_));
 sky130_fd_sc_hd__mux2_1 _7423_ (.A0(\ann.ReLU_out[9][13] ),
    .A1(_3763_),
    .S(net39),
    .X(_3764_));
 sky130_fd_sc_hd__mux2_1 _7424_ (.A0(net315),
    .A1(_3764_),
    .S(net89),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _7425_ (.A0(\ann.ReLU_out[1][14] ),
    .A1(\ann.ReLU_out[0][14] ),
    .S(net40),
    .X(_3765_));
 sky130_fd_sc_hd__mux2_1 _7426_ (.A0(\ann.ReLU_out[2][14] ),
    .A1(_3765_),
    .S(net42),
    .X(_3766_));
 sky130_fd_sc_hd__mux2_1 _7427_ (.A0(\ann.ReLU_out[3][14] ),
    .A1(_3766_),
    .S(net36),
    .X(_3767_));
 sky130_fd_sc_hd__mux2_1 _7428_ (.A0(_3767_),
    .A1(\ann.ReLU_out[4][14] ),
    .S(net54),
    .X(_3768_));
 sky130_fd_sc_hd__mux2_1 _7429_ (.A0(_3768_),
    .A1(\ann.ReLU_out[5][14] ),
    .S(net56),
    .X(_3769_));
 sky130_fd_sc_hd__mux2_1 _7430_ (.A0(_3769_),
    .A1(\ann.ReLU_out[6][14] ),
    .S(net45),
    .X(_3770_));
 sky130_fd_sc_hd__mux2_1 _7431_ (.A0(_3770_),
    .A1(\ann.ReLU_out[7][14] ),
    .S(net48),
    .X(_3771_));
 sky130_fd_sc_hd__mux2_1 _7432_ (.A0(\ann.ReLU_out[8][14] ),
    .A1(_3771_),
    .S(net51),
    .X(_3772_));
 sky130_fd_sc_hd__mux2_1 _7433_ (.A0(\ann.ReLU_out[9][14] ),
    .A1(_3772_),
    .S(net39),
    .X(_3773_));
 sky130_fd_sc_hd__mux2_1 _7434_ (.A0(net313),
    .A1(_3773_),
    .S(net89),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _7435_ (.A0(\ann.ReLU_out[1][15] ),
    .A1(\ann.ReLU_out[0][15] ),
    .S(net40),
    .X(_3774_));
 sky130_fd_sc_hd__mux2_1 _7436_ (.A0(\ann.ReLU_out[2][15] ),
    .A1(_3774_),
    .S(net42),
    .X(_3775_));
 sky130_fd_sc_hd__mux2_1 _7437_ (.A0(\ann.ReLU_out[3][15] ),
    .A1(_3775_),
    .S(net36),
    .X(_3776_));
 sky130_fd_sc_hd__mux2_1 _7438_ (.A0(_3776_),
    .A1(\ann.ReLU_out[4][15] ),
    .S(net54),
    .X(_3777_));
 sky130_fd_sc_hd__mux2_1 _7439_ (.A0(_3777_),
    .A1(\ann.ReLU_out[5][15] ),
    .S(net56),
    .X(_3778_));
 sky130_fd_sc_hd__mux2_1 _7440_ (.A0(_3778_),
    .A1(net677),
    .S(net45),
    .X(_3779_));
 sky130_fd_sc_hd__mux2_1 _7441_ (.A0(_3779_),
    .A1(net687),
    .S(net48),
    .X(_3780_));
 sky130_fd_sc_hd__mux2_1 _7442_ (.A0(net669),
    .A1(_3780_),
    .S(net51),
    .X(_3781_));
 sky130_fd_sc_hd__mux2_1 _7443_ (.A0(net682),
    .A1(_3781_),
    .S(net39),
    .X(_3782_));
 sky130_fd_sc_hd__mux2_1 _7444_ (.A0(net712),
    .A1(_3782_),
    .S(net89),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _7445_ (.A0(\ann.ReLU_out[1][16] ),
    .A1(\ann.ReLU_out[0][16] ),
    .S(net40),
    .X(_3783_));
 sky130_fd_sc_hd__mux2_1 _7446_ (.A0(\ann.ReLU_out[2][16] ),
    .A1(_3783_),
    .S(net42),
    .X(_3784_));
 sky130_fd_sc_hd__mux2_1 _7447_ (.A0(\ann.ReLU_out[3][16] ),
    .A1(_3784_),
    .S(net36),
    .X(_3785_));
 sky130_fd_sc_hd__mux2_1 _7448_ (.A0(_3785_),
    .A1(net412),
    .S(net53),
    .X(_3786_));
 sky130_fd_sc_hd__mux2_1 _7449_ (.A0(_3786_),
    .A1(net440),
    .S(net55),
    .X(_3787_));
 sky130_fd_sc_hd__a21oi_1 _7450_ (.A1(_0680_),
    .A2(net44),
    .B1(net47),
    .Y(_3788_));
 sky130_fd_sc_hd__o21a_1 _7451_ (.A1(net44),
    .A2(_3787_),
    .B1(_3788_),
    .X(_3789_));
 sky130_fd_sc_hd__a21bo_1 _7452_ (.A1(net538),
    .A2(net47),
    .B1_N(net50),
    .X(_3790_));
 sky130_fd_sc_hd__o22a_1 _7453_ (.A1(net464),
    .A2(net50),
    .B1(_3789_),
    .B2(_3790_),
    .X(_3791_));
 sky130_fd_sc_hd__mux2_1 _7454_ (.A0(net452),
    .A1(_3791_),
    .S(net38),
    .X(_3792_));
 sky130_fd_sc_hd__mux2_1 _7455_ (.A0(net755),
    .A1(_3792_),
    .S(net89),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _7456_ (.A0(\ann.ReLU_out[1][17] ),
    .A1(\ann.ReLU_out[0][17] ),
    .S(net40),
    .X(_3793_));
 sky130_fd_sc_hd__mux2_1 _7457_ (.A0(\ann.ReLU_out[2][17] ),
    .A1(_3793_),
    .S(net43),
    .X(_3794_));
 sky130_fd_sc_hd__mux2_1 _7458_ (.A0(\ann.ReLU_out[3][17] ),
    .A1(_3794_),
    .S(net37),
    .X(_3795_));
 sky130_fd_sc_hd__mux2_1 _7459_ (.A0(_3795_),
    .A1(net439),
    .S(net54),
    .X(_3796_));
 sky130_fd_sc_hd__mux2_1 _7460_ (.A0(_3796_),
    .A1(net527),
    .S(net55),
    .X(_3797_));
 sky130_fd_sc_hd__a21oi_1 _7461_ (.A1(_0679_),
    .A2(net44),
    .B1(net48),
    .Y(_3798_));
 sky130_fd_sc_hd__o21a_1 _7462_ (.A1(net44),
    .A2(_3797_),
    .B1(_3798_),
    .X(_3799_));
 sky130_fd_sc_hd__a21bo_1 _7463_ (.A1(net637),
    .A2(net47),
    .B1_N(net50),
    .X(_3800_));
 sky130_fd_sc_hd__o22a_1 _7464_ (.A1(net587),
    .A2(net50),
    .B1(_3799_),
    .B2(_3800_),
    .X(_3801_));
 sky130_fd_sc_hd__mux2_1 _7465_ (.A0(net406),
    .A1(_3801_),
    .S(net38),
    .X(_3802_));
 sky130_fd_sc_hd__mux2_1 _7466_ (.A0(net188),
    .A1(_3802_),
    .S(net90),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _7467_ (.A0(\ann.ReLU_out[1][18] ),
    .A1(\ann.ReLU_out[0][18] ),
    .S(net41),
    .X(_3803_));
 sky130_fd_sc_hd__mux2_1 _7468_ (.A0(\ann.ReLU_out[2][18] ),
    .A1(_3803_),
    .S(net43),
    .X(_3804_));
 sky130_fd_sc_hd__mux2_1 _7469_ (.A0(\ann.ReLU_out[3][18] ),
    .A1(_3804_),
    .S(net36),
    .X(_3805_));
 sky130_fd_sc_hd__mux2_1 _7470_ (.A0(_3805_),
    .A1(\ann.ReLU_out[4][18] ),
    .S(net53),
    .X(_3806_));
 sky130_fd_sc_hd__mux2_1 _7471_ (.A0(_3806_),
    .A1(\ann.ReLU_out[5][18] ),
    .S(net55),
    .X(_3807_));
 sky130_fd_sc_hd__mux2_1 _7472_ (.A0(_3807_),
    .A1(net463),
    .S(net44),
    .X(_3808_));
 sky130_fd_sc_hd__mux2_1 _7473_ (.A0(_3808_),
    .A1(net679),
    .S(net47),
    .X(_3809_));
 sky130_fd_sc_hd__mux2_1 _7474_ (.A0(net708),
    .A1(_3809_),
    .S(net50),
    .X(_3810_));
 sky130_fd_sc_hd__mux2_1 _7475_ (.A0(net636),
    .A1(_3810_),
    .S(net38),
    .X(_3811_));
 sky130_fd_sc_hd__mux2_1 _7476_ (.A0(net187),
    .A1(_3811_),
    .S(net90),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _7477_ (.A0(\ann.ReLU_out[1][19] ),
    .A1(\ann.ReLU_out[0][19] ),
    .S(net40),
    .X(_3812_));
 sky130_fd_sc_hd__mux2_1 _7478_ (.A0(\ann.ReLU_out[2][19] ),
    .A1(_3812_),
    .S(net42),
    .X(_3813_));
 sky130_fd_sc_hd__mux2_1 _7479_ (.A0(\ann.ReLU_out[3][19] ),
    .A1(_3813_),
    .S(net36),
    .X(_3814_));
 sky130_fd_sc_hd__mux2_1 _7480_ (.A0(_3814_),
    .A1(\ann.ReLU_out[4][19] ),
    .S(net53),
    .X(_3815_));
 sky130_fd_sc_hd__mux2_1 _7481_ (.A0(_3815_),
    .A1(\ann.ReLU_out[5][19] ),
    .S(net55),
    .X(_3816_));
 sky130_fd_sc_hd__mux2_1 _7482_ (.A0(_3816_),
    .A1(net655),
    .S(net44),
    .X(_3817_));
 sky130_fd_sc_hd__mux2_1 _7483_ (.A0(_3817_),
    .A1(net641),
    .S(net47),
    .X(_3818_));
 sky130_fd_sc_hd__mux2_1 _7484_ (.A0(net646),
    .A1(_3818_),
    .S(net50),
    .X(_3819_));
 sky130_fd_sc_hd__mux2_1 _7485_ (.A0(net673),
    .A1(_3819_),
    .S(net38),
    .X(_3820_));
 sky130_fd_sc_hd__mux2_1 _7486_ (.A0(net774),
    .A1(_3820_),
    .S(net89),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _7487_ (.A0(\ann.ReLU_out[1][20] ),
    .A1(\ann.ReLU_out[0][20] ),
    .S(_3629_),
    .X(_3821_));
 sky130_fd_sc_hd__mux2_1 _7488_ (.A0(\ann.ReLU_out[2][20] ),
    .A1(_3821_),
    .S(_3566_),
    .X(_3822_));
 sky130_fd_sc_hd__mux2_1 _7489_ (.A0(\ann.ReLU_out[3][20] ),
    .A1(_3822_),
    .S(_3507_),
    .X(_3823_));
 sky130_fd_sc_hd__mux2_1 _7490_ (.A0(_3823_),
    .A1(\ann.ReLU_out[4][20] ),
    .S(net53),
    .X(_3824_));
 sky130_fd_sc_hd__mux2_1 _7491_ (.A0(_3824_),
    .A1(\ann.ReLU_out[5][20] ),
    .S(net55),
    .X(_3825_));
 sky130_fd_sc_hd__mux2_1 _7492_ (.A0(_3825_),
    .A1(net651),
    .S(net44),
    .X(_3826_));
 sky130_fd_sc_hd__mux2_1 _7493_ (.A0(_3826_),
    .A1(net663),
    .S(net47),
    .X(_3827_));
 sky130_fd_sc_hd__mux2_1 _7494_ (.A0(net634),
    .A1(_3827_),
    .S(net50),
    .X(_3828_));
 sky130_fd_sc_hd__mux2_1 _7495_ (.A0(net659),
    .A1(_3828_),
    .S(net38),
    .X(_3829_));
 sky130_fd_sc_hd__mux2_1 _7496_ (.A0(net666),
    .A1(_3829_),
    .S(net89),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _7497_ (.A0(\ann.ReLU_out[1][21] ),
    .A1(\ann.ReLU_out[0][21] ),
    .S(net41),
    .X(_3830_));
 sky130_fd_sc_hd__mux2_1 _7498_ (.A0(\ann.ReLU_out[2][21] ),
    .A1(_3830_),
    .S(net43),
    .X(_3831_));
 sky130_fd_sc_hd__mux2_1 _7499_ (.A0(\ann.ReLU_out[3][21] ),
    .A1(_3831_),
    .S(net37),
    .X(_3832_));
 sky130_fd_sc_hd__mux2_1 _7500_ (.A0(_3832_),
    .A1(\ann.ReLU_out[4][21] ),
    .S(net53),
    .X(_3833_));
 sky130_fd_sc_hd__mux2_1 _7501_ (.A0(_3833_),
    .A1(\ann.ReLU_out[5][21] ),
    .S(net55),
    .X(_3834_));
 sky130_fd_sc_hd__mux2_1 _7502_ (.A0(_3834_),
    .A1(net475),
    .S(net44),
    .X(_3835_));
 sky130_fd_sc_hd__mux2_1 _7503_ (.A0(_3835_),
    .A1(net633),
    .S(net47),
    .X(_3836_));
 sky130_fd_sc_hd__mux2_1 _7504_ (.A0(net632),
    .A1(_3836_),
    .S(net50),
    .X(_3837_));
 sky130_fd_sc_hd__mux2_1 _7505_ (.A0(net599),
    .A1(_3837_),
    .S(net38),
    .X(_3838_));
 sky130_fd_sc_hd__mux2_1 _7506_ (.A0(net675),
    .A1(_3838_),
    .S(net89),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _7507_ (.A0(\ann.ReLU_out[1][22] ),
    .A1(\ann.ReLU_out[0][22] ),
    .S(net41),
    .X(_3839_));
 sky130_fd_sc_hd__mux2_1 _7508_ (.A0(\ann.ReLU_out[2][22] ),
    .A1(_3839_),
    .S(net43),
    .X(_3840_));
 sky130_fd_sc_hd__mux2_1 _7509_ (.A0(\ann.ReLU_out[3][22] ),
    .A1(_3840_),
    .S(net37),
    .X(_3841_));
 sky130_fd_sc_hd__mux2_1 _7510_ (.A0(_3841_),
    .A1(\ann.ReLU_out[4][22] ),
    .S(net54),
    .X(_3842_));
 sky130_fd_sc_hd__mux2_1 _7511_ (.A0(_3842_),
    .A1(net422),
    .S(net55),
    .X(_3843_));
 sky130_fd_sc_hd__mux2_1 _7512_ (.A0(_3843_),
    .A1(net399),
    .S(net44),
    .X(_3844_));
 sky130_fd_sc_hd__mux2_1 _7513_ (.A0(_3844_),
    .A1(net483),
    .S(net47),
    .X(_3845_));
 sky130_fd_sc_hd__mux2_1 _7514_ (.A0(net478),
    .A1(_3845_),
    .S(net50),
    .X(_3846_));
 sky130_fd_sc_hd__mux2_1 _7515_ (.A0(net657),
    .A1(_3846_),
    .S(net38),
    .X(_3847_));
 sky130_fd_sc_hd__mux2_1 _7516_ (.A0(net186),
    .A1(_3847_),
    .S(net90),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _7517_ (.A0(\ann.ReLU_out[1][23] ),
    .A1(\ann.ReLU_out[0][23] ),
    .S(net41),
    .X(_3848_));
 sky130_fd_sc_hd__mux2_1 _7518_ (.A0(\ann.ReLU_out[2][23] ),
    .A1(_3848_),
    .S(net43),
    .X(_3849_));
 sky130_fd_sc_hd__mux2_1 _7519_ (.A0(\ann.ReLU_out[3][23] ),
    .A1(_3849_),
    .S(net37),
    .X(_3850_));
 sky130_fd_sc_hd__mux2_1 _7520_ (.A0(_3850_),
    .A1(\ann.ReLU_out[4][23] ),
    .S(net54),
    .X(_3851_));
 sky130_fd_sc_hd__mux2_1 _7521_ (.A0(_3851_),
    .A1(\ann.ReLU_out[5][23] ),
    .S(net56),
    .X(_3852_));
 sky130_fd_sc_hd__mux2_1 _7522_ (.A0(_3852_),
    .A1(net493),
    .S(net46),
    .X(_3853_));
 sky130_fd_sc_hd__mux2_1 _7523_ (.A0(_3853_),
    .A1(net424),
    .S(net49),
    .X(_3854_));
 sky130_fd_sc_hd__mux2_1 _7524_ (.A0(net418),
    .A1(_3854_),
    .S(net52),
    .X(_3855_));
 sky130_fd_sc_hd__mux2_1 _7525_ (.A0(net453),
    .A1(_3855_),
    .S(net39),
    .X(_3856_));
 sky130_fd_sc_hd__mux2_1 _7526_ (.A0(net658),
    .A1(_3856_),
    .S(net90),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _7527_ (.A0(\ann.ReLU_out[1][24] ),
    .A1(\ann.ReLU_out[0][24] ),
    .S(net41),
    .X(_3857_));
 sky130_fd_sc_hd__mux2_1 _7528_ (.A0(\ann.ReLU_out[2][24] ),
    .A1(_3857_),
    .S(net43),
    .X(_3858_));
 sky130_fd_sc_hd__mux2_1 _7529_ (.A0(\ann.ReLU_out[3][24] ),
    .A1(_3858_),
    .S(net37),
    .X(_3859_));
 sky130_fd_sc_hd__mux2_1 _7530_ (.A0(_3859_),
    .A1(\ann.ReLU_out[4][24] ),
    .S(net54),
    .X(_3860_));
 sky130_fd_sc_hd__mux2_1 _7531_ (.A0(_3860_),
    .A1(net447),
    .S(net56),
    .X(_3861_));
 sky130_fd_sc_hd__mux2_1 _7532_ (.A0(_3861_),
    .A1(net446),
    .S(net46),
    .X(_3862_));
 sky130_fd_sc_hd__mux2_1 _7533_ (.A0(_3862_),
    .A1(net428),
    .S(net49),
    .X(_3863_));
 sky130_fd_sc_hd__mux2_1 _7534_ (.A0(net411),
    .A1(_3863_),
    .S(net52),
    .X(_3864_));
 sky130_fd_sc_hd__mux2_1 _7535_ (.A0(net548),
    .A1(_3864_),
    .S(net39),
    .X(_3865_));
 sky130_fd_sc_hd__mux2_1 _7536_ (.A0(net644),
    .A1(_3865_),
    .S(net90),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _7537_ (.A0(\ann.ReLU_out[1][25] ),
    .A1(\ann.ReLU_out[0][25] ),
    .S(net41),
    .X(_3866_));
 sky130_fd_sc_hd__mux2_1 _7538_ (.A0(\ann.ReLU_out[2][25] ),
    .A1(_3866_),
    .S(net43),
    .X(_3867_));
 sky130_fd_sc_hd__mux2_1 _7539_ (.A0(\ann.ReLU_out[3][25] ),
    .A1(_3867_),
    .S(net37),
    .X(_3868_));
 sky130_fd_sc_hd__mux2_1 _7540_ (.A0(_3868_),
    .A1(\ann.ReLU_out[4][25] ),
    .S(net53),
    .X(_3869_));
 sky130_fd_sc_hd__mux2_1 _7541_ (.A0(_3869_),
    .A1(\ann.ReLU_out[5][25] ),
    .S(net55),
    .X(_3870_));
 sky130_fd_sc_hd__mux2_1 _7542_ (.A0(_3870_),
    .A1(net529),
    .S(net46),
    .X(_3871_));
 sky130_fd_sc_hd__mux2_1 _7543_ (.A0(_3871_),
    .A1(net425),
    .S(net49),
    .X(_3872_));
 sky130_fd_sc_hd__mux2_1 _7544_ (.A0(net517),
    .A1(_3872_),
    .S(net52),
    .X(_3873_));
 sky130_fd_sc_hd__mux2_1 _7545_ (.A0(net608),
    .A1(_3873_),
    .S(net39),
    .X(_3874_));
 sky130_fd_sc_hd__mux2_1 _7546_ (.A0(net656),
    .A1(_3874_),
    .S(net90),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _7547_ (.A0(\ann.ReLU_out[1][26] ),
    .A1(\ann.ReLU_out[0][26] ),
    .S(net40),
    .X(_3875_));
 sky130_fd_sc_hd__mux2_1 _7548_ (.A0(\ann.ReLU_out[2][26] ),
    .A1(_3875_),
    .S(net42),
    .X(_3876_));
 sky130_fd_sc_hd__mux2_1 _7549_ (.A0(\ann.ReLU_out[3][26] ),
    .A1(_3876_),
    .S(net37),
    .X(_3877_));
 sky130_fd_sc_hd__mux2_1 _7550_ (.A0(_3877_),
    .A1(\ann.ReLU_out[4][26] ),
    .S(_3444_),
    .X(_3878_));
 sky130_fd_sc_hd__mux2_1 _7551_ (.A0(_3878_),
    .A1(net534),
    .S(net55),
    .X(_3879_));
 sky130_fd_sc_hd__mux2_1 _7552_ (.A0(_3879_),
    .A1(net487),
    .S(net46),
    .X(_3880_));
 sky130_fd_sc_hd__mux2_1 _7553_ (.A0(_3880_),
    .A1(net501),
    .S(net47),
    .X(_3881_));
 sky130_fd_sc_hd__mux2_1 _7554_ (.A0(net455),
    .A1(_3881_),
    .S(net52),
    .X(_3882_));
 sky130_fd_sc_hd__mux2_1 _7555_ (.A0(net581),
    .A1(_3882_),
    .S(net39),
    .X(_3883_));
 sky130_fd_sc_hd__mux2_1 _7556_ (.A0(net182),
    .A1(_3883_),
    .S(net90),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _7557_ (.A0(\ann.ReLU_out[1][27] ),
    .A1(\ann.ReLU_out[0][27] ),
    .S(net40),
    .X(_3884_));
 sky130_fd_sc_hd__mux2_1 _7558_ (.A0(\ann.ReLU_out[2][27] ),
    .A1(_3884_),
    .S(net42),
    .X(_3885_));
 sky130_fd_sc_hd__mux2_1 _7559_ (.A0(\ann.ReLU_out[3][27] ),
    .A1(_3885_),
    .S(net36),
    .X(_3886_));
 sky130_fd_sc_hd__mux2_1 _7560_ (.A0(_3886_),
    .A1(\ann.ReLU_out[4][27] ),
    .S(net53),
    .X(_3887_));
 sky130_fd_sc_hd__mux2_1 _7561_ (.A0(_3887_),
    .A1(net624),
    .S(net55),
    .X(_3888_));
 sky130_fd_sc_hd__mux2_1 _7562_ (.A0(_3888_),
    .A1(net481),
    .S(net46),
    .X(_3889_));
 sky130_fd_sc_hd__mux2_1 _7563_ (.A0(_3889_),
    .A1(net627),
    .S(net47),
    .X(_3890_));
 sky130_fd_sc_hd__mux2_1 _7564_ (.A0(net643),
    .A1(_3890_),
    .S(net50),
    .X(_3891_));
 sky130_fd_sc_hd__mux2_1 _7565_ (.A0(net664),
    .A1(_3891_),
    .S(net38),
    .X(_3892_));
 sky130_fd_sc_hd__mux2_1 _7566_ (.A0(net757),
    .A1(_3892_),
    .S(_3637_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _7567_ (.A0(\ann.ReLU_out[1][28] ),
    .A1(\ann.ReLU_out[0][28] ),
    .S(net40),
    .X(_3893_));
 sky130_fd_sc_hd__mux2_1 _7568_ (.A0(\ann.ReLU_out[2][28] ),
    .A1(_3893_),
    .S(net42),
    .X(_3894_));
 sky130_fd_sc_hd__mux2_1 _7569_ (.A0(\ann.ReLU_out[3][28] ),
    .A1(_3894_),
    .S(net36),
    .X(_3895_));
 sky130_fd_sc_hd__mux2_1 _7570_ (.A0(_3895_),
    .A1(\ann.ReLU_out[4][28] ),
    .S(net53),
    .X(_3896_));
 sky130_fd_sc_hd__mux2_1 _7571_ (.A0(_3896_),
    .A1(net609),
    .S(net55),
    .X(_3897_));
 sky130_fd_sc_hd__mux2_1 _7572_ (.A0(_3897_),
    .A1(net568),
    .S(net44),
    .X(_3898_));
 sky130_fd_sc_hd__mux2_1 _7573_ (.A0(_3898_),
    .A1(net593),
    .S(net47),
    .X(_3899_));
 sky130_fd_sc_hd__mux2_1 _7574_ (.A0(net586),
    .A1(_3899_),
    .S(net50),
    .X(_3900_));
 sky130_fd_sc_hd__mux2_1 _7575_ (.A0(net462),
    .A1(_3900_),
    .S(net38),
    .X(_3901_));
 sky130_fd_sc_hd__mux2_1 _7576_ (.A0(net743),
    .A1(_3901_),
    .S(net89),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _7577_ (.A0(\ann.ReLU_out[1][29] ),
    .A1(\ann.ReLU_out[0][29] ),
    .S(net40),
    .X(_3902_));
 sky130_fd_sc_hd__mux2_1 _7578_ (.A0(\ann.ReLU_out[2][29] ),
    .A1(_3902_),
    .S(net42),
    .X(_3903_));
 sky130_fd_sc_hd__mux2_1 _7579_ (.A0(\ann.ReLU_out[3][29] ),
    .A1(_3903_),
    .S(net36),
    .X(_3904_));
 sky130_fd_sc_hd__mux2_1 _7580_ (.A0(_3904_),
    .A1(\ann.ReLU_out[4][29] ),
    .S(net53),
    .X(_3905_));
 sky130_fd_sc_hd__mux2_1 _7581_ (.A0(_3905_),
    .A1(\ann.ReLU_out[5][29] ),
    .S(net55),
    .X(_3906_));
 sky130_fd_sc_hd__mux2_1 _7582_ (.A0(_3906_),
    .A1(net498),
    .S(net44),
    .X(_3907_));
 sky130_fd_sc_hd__mux2_1 _7583_ (.A0(_3907_),
    .A1(net640),
    .S(net47),
    .X(_3908_));
 sky130_fd_sc_hd__mux2_1 _7584_ (.A0(net676),
    .A1(_3908_),
    .S(net50),
    .X(_3909_));
 sky130_fd_sc_hd__mux2_1 _7585_ (.A0(net672),
    .A1(_3909_),
    .S(net38),
    .X(_3910_));
 sky130_fd_sc_hd__mux2_1 _7586_ (.A0(net717),
    .A1(_3910_),
    .S(net89),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _7587_ (.A0(\ann.ReLU_out[1][30] ),
    .A1(\ann.ReLU_out[0][30] ),
    .S(net40),
    .X(_3911_));
 sky130_fd_sc_hd__mux2_1 _7588_ (.A0(\ann.ReLU_out[2][30] ),
    .A1(_3911_),
    .S(net42),
    .X(_3912_));
 sky130_fd_sc_hd__mux2_1 _7589_ (.A0(\ann.ReLU_out[3][30] ),
    .A1(_3912_),
    .S(net36),
    .X(_3913_));
 sky130_fd_sc_hd__mux2_1 _7590_ (.A0(_3913_),
    .A1(\ann.ReLU_out[4][30] ),
    .S(net53),
    .X(_3914_));
 sky130_fd_sc_hd__mux2_1 _7591_ (.A0(_3914_),
    .A1(\ann.ReLU_out[5][30] ),
    .S(net55),
    .X(_3915_));
 sky130_fd_sc_hd__or2_1 _7592_ (.A(net44),
    .B(_3915_),
    .X(_3916_));
 sky130_fd_sc_hd__a21oi_1 _7593_ (.A1(_0597_),
    .A2(net44),
    .B1(net47),
    .Y(_3917_));
 sky130_fd_sc_hd__a22o_1 _7594_ (.A1(net613),
    .A2(net47),
    .B1(_3916_),
    .B2(_3917_),
    .X(_3918_));
 sky130_fd_sc_hd__mux2_1 _7595_ (.A0(net610),
    .A1(_3918_),
    .S(net50),
    .X(_3919_));
 sky130_fd_sc_hd__inv_2 _7596_ (.A(_3919_),
    .Y(_3920_));
 sky130_fd_sc_hd__o21ai_1 _7597_ (.A1(net631),
    .A2(net38),
    .B1(net89),
    .Y(_3921_));
 sky130_fd_sc_hd__a21o_1 _7598_ (.A1(net38),
    .A2(_3920_),
    .B1(_3921_),
    .X(_3922_));
 sky130_fd_sc_hd__o21ai_1 _7599_ (.A1(net104),
    .A2(net89),
    .B1(_3922_),
    .Y(_0134_));
 sky130_fd_sc_hd__nor2_1 _7600_ (.A(net18),
    .B(net17),
    .Y(_3923_));
 sky130_fd_sc_hd__a41o_1 _7601_ (.A1(_0560_),
    .A2(_0561_),
    .A3(net20),
    .A4(_3923_),
    .B1(net31),
    .X(_3924_));
 sky130_fd_sc_hd__and2b_2 _7602_ (.A_N(net58),
    .B(\ann.sum[0] ),
    .X(_3925_));
 sky130_fd_sc_hd__mux2_1 _7603_ (.A0(net287),
    .A1(_3925_),
    .S(net88),
    .X(_0135_));
 sky130_fd_sc_hd__and2b_2 _7604_ (.A_N(net58),
    .B(\ann.sum[1] ),
    .X(_3926_));
 sky130_fd_sc_hd__mux2_1 _7605_ (.A0(net263),
    .A1(_3926_),
    .S(net88),
    .X(_0136_));
 sky130_fd_sc_hd__and2b_2 _7606_ (.A_N(net58),
    .B(\ann.sum[2] ),
    .X(_3927_));
 sky130_fd_sc_hd__mux2_1 _7607_ (.A0(net283),
    .A1(_3927_),
    .S(net88),
    .X(_0137_));
 sky130_fd_sc_hd__and2b_2 _7608_ (.A_N(net58),
    .B(\ann.sum[3] ),
    .X(_3928_));
 sky130_fd_sc_hd__mux2_1 _7609_ (.A0(net303),
    .A1(_3928_),
    .S(net88),
    .X(_0138_));
 sky130_fd_sc_hd__and2b_2 _7610_ (.A_N(net58),
    .B(\ann.sum[4] ),
    .X(_3929_));
 sky130_fd_sc_hd__mux2_1 _7611_ (.A0(net295),
    .A1(_3929_),
    .S(net88),
    .X(_0139_));
 sky130_fd_sc_hd__and2b_2 _7612_ (.A_N(net58),
    .B(\ann.sum[5] ),
    .X(_3930_));
 sky130_fd_sc_hd__mux2_1 _7613_ (.A0(net297),
    .A1(_3930_),
    .S(net88),
    .X(_0140_));
 sky130_fd_sc_hd__and2b_2 _7614_ (.A_N(net58),
    .B(\ann.sum[6] ),
    .X(_3931_));
 sky130_fd_sc_hd__mux2_1 _7615_ (.A0(net291),
    .A1(_3931_),
    .S(net88),
    .X(_0141_));
 sky130_fd_sc_hd__and2b_4 _7616_ (.A_N(net59),
    .B(\ann.sum[7] ),
    .X(_3932_));
 sky130_fd_sc_hd__mux2_1 _7617_ (.A0(net277),
    .A1(_3932_),
    .S(net88),
    .X(_0142_));
 sky130_fd_sc_hd__and2b_4 _7618_ (.A_N(net58),
    .B(\ann.sum[8] ),
    .X(_3933_));
 sky130_fd_sc_hd__mux2_1 _7619_ (.A0(net305),
    .A1(_3933_),
    .S(net87),
    .X(_0143_));
 sky130_fd_sc_hd__and2b_4 _7620_ (.A_N(net58),
    .B(\ann.sum[9] ),
    .X(_3934_));
 sky130_fd_sc_hd__mux2_1 _7621_ (.A0(net261),
    .A1(_3934_),
    .S(net87),
    .X(_0144_));
 sky130_fd_sc_hd__and2b_4 _7622_ (.A_N(net58),
    .B(\ann.sum[10] ),
    .X(_3935_));
 sky130_fd_sc_hd__mux2_1 _7623_ (.A0(net275),
    .A1(_3935_),
    .S(net87),
    .X(_0145_));
 sky130_fd_sc_hd__and2b_4 _7624_ (.A_N(\ann.sum[31] ),
    .B(\ann.sum[11] ),
    .X(_3936_));
 sky130_fd_sc_hd__mux2_1 _7625_ (.A0(net301),
    .A1(_3936_),
    .S(net87),
    .X(_0146_));
 sky130_fd_sc_hd__and2b_4 _7626_ (.A_N(\ann.sum[31] ),
    .B(\ann.sum[12] ),
    .X(_3937_));
 sky130_fd_sc_hd__mux2_1 _7627_ (.A0(net269),
    .A1(_3937_),
    .S(net87),
    .X(_0147_));
 sky130_fd_sc_hd__and2b_4 _7628_ (.A_N(net58),
    .B(\ann.sum[13] ),
    .X(_3938_));
 sky130_fd_sc_hd__mux2_1 _7629_ (.A0(net265),
    .A1(_3938_),
    .S(net87),
    .X(_0148_));
 sky130_fd_sc_hd__and2b_4 _7630_ (.A_N(net58),
    .B(\ann.sum[14] ),
    .X(_3939_));
 sky130_fd_sc_hd__mux2_1 _7631_ (.A0(net259),
    .A1(_3939_),
    .S(net88),
    .X(_0149_));
 sky130_fd_sc_hd__and2b_4 _7632_ (.A_N(net58),
    .B(\ann.sum[15] ),
    .X(_3940_));
 sky130_fd_sc_hd__mux2_1 _7633_ (.A0(net317),
    .A1(_3940_),
    .S(net87),
    .X(_0150_));
 sky130_fd_sc_hd__and2b_4 _7634_ (.A_N(net58),
    .B(\ann.sum[16] ),
    .X(_3941_));
 sky130_fd_sc_hd__mux2_1 _7635_ (.A0(net279),
    .A1(_3941_),
    .S(net87),
    .X(_0151_));
 sky130_fd_sc_hd__and2b_4 _7636_ (.A_N(net58),
    .B(\ann.sum[17] ),
    .X(_3942_));
 sky130_fd_sc_hd__mux2_1 _7637_ (.A0(net271),
    .A1(_3942_),
    .S(net87),
    .X(_0152_));
 sky130_fd_sc_hd__and2b_4 _7638_ (.A_N(net58),
    .B(\ann.sum[18] ),
    .X(_3943_));
 sky130_fd_sc_hd__mux2_1 _7639_ (.A0(net267),
    .A1(_3943_),
    .S(net87),
    .X(_0153_));
 sky130_fd_sc_hd__and2b_4 _7640_ (.A_N(net59),
    .B(\ann.sum[19] ),
    .X(_3944_));
 sky130_fd_sc_hd__mux2_1 _7641_ (.A0(net307),
    .A1(_3944_),
    .S(net87),
    .X(_0154_));
 sky130_fd_sc_hd__and2b_4 _7642_ (.A_N(net59),
    .B(\ann.sum[20] ),
    .X(_3945_));
 sky130_fd_sc_hd__mux2_1 _7643_ (.A0(net285),
    .A1(_3945_),
    .S(net88),
    .X(_0155_));
 sky130_fd_sc_hd__and2b_4 _7644_ (.A_N(net59),
    .B(\ann.sum[21] ),
    .X(_3946_));
 sky130_fd_sc_hd__mux2_1 _7645_ (.A0(net255),
    .A1(_3946_),
    .S(net88),
    .X(_0156_));
 sky130_fd_sc_hd__and2b_4 _7646_ (.A_N(net59),
    .B(\ann.sum[22] ),
    .X(_3947_));
 sky130_fd_sc_hd__mux2_1 _7647_ (.A0(net299),
    .A1(_3947_),
    .S(net88),
    .X(_0157_));
 sky130_fd_sc_hd__and2b_4 _7648_ (.A_N(net59),
    .B(\ann.sum[23] ),
    .X(_3948_));
 sky130_fd_sc_hd__mux2_1 _7649_ (.A0(net281),
    .A1(_3948_),
    .S(net88),
    .X(_0158_));
 sky130_fd_sc_hd__and2b_2 _7650_ (.A_N(net59),
    .B(\ann.sum[24] ),
    .X(_3949_));
 sky130_fd_sc_hd__mux2_1 _7651_ (.A0(net289),
    .A1(_3949_),
    .S(net88),
    .X(_0159_));
 sky130_fd_sc_hd__and2b_4 _7652_ (.A_N(net59),
    .B(\ann.sum[25] ),
    .X(_3950_));
 sky130_fd_sc_hd__mux2_1 _7653_ (.A0(net309),
    .A1(_3950_),
    .S(net88),
    .X(_0160_));
 sky130_fd_sc_hd__and2b_4 _7654_ (.A_N(net59),
    .B(\ann.sum[26] ),
    .X(_3951_));
 sky130_fd_sc_hd__mux2_1 _7655_ (.A0(net319),
    .A1(_3951_),
    .S(net87),
    .X(_0161_));
 sky130_fd_sc_hd__and2b_4 _7656_ (.A_N(net59),
    .B(\ann.sum[27] ),
    .X(_3952_));
 sky130_fd_sc_hd__mux2_1 _7657_ (.A0(net293),
    .A1(_3952_),
    .S(net87),
    .X(_0162_));
 sky130_fd_sc_hd__and2b_4 _7658_ (.A_N(net59),
    .B(\ann.sum[28] ),
    .X(_3953_));
 sky130_fd_sc_hd__mux2_1 _7659_ (.A0(net311),
    .A1(_3953_),
    .S(net87),
    .X(_0163_));
 sky130_fd_sc_hd__and2b_4 _7660_ (.A_N(net59),
    .B(\ann.sum[29] ),
    .X(_3954_));
 sky130_fd_sc_hd__mux2_1 _7661_ (.A0(net273),
    .A1(_3954_),
    .S(net87),
    .X(_0164_));
 sky130_fd_sc_hd__and2b_4 _7662_ (.A_N(net59),
    .B(\ann.sum[30] ),
    .X(_3955_));
 sky130_fd_sc_hd__mux2_1 _7663_ (.A0(net257),
    .A1(_3955_),
    .S(net87),
    .X(_0165_));
 sky130_fd_sc_hd__a41o_1 _7664_ (.A1(_0560_),
    .A2(net15),
    .A3(net20),
    .A4(_3923_),
    .B1(net31),
    .X(_3956_));
 sky130_fd_sc_hd__mux2_1 _7665_ (.A0(net323),
    .A1(_3925_),
    .S(net86),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _7666_ (.A0(net573),
    .A1(_3926_),
    .S(net86),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _7667_ (.A0(net520),
    .A1(_3927_),
    .S(net86),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _7668_ (.A0(net540),
    .A1(_3928_),
    .S(net86),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _7669_ (.A0(net566),
    .A1(_3929_),
    .S(net86),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _7670_ (.A0(net537),
    .A1(_3930_),
    .S(net86),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _7671_ (.A0(net522),
    .A1(_3931_),
    .S(net86),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _7672_ (.A0(net561),
    .A1(_3932_),
    .S(net86),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _7673_ (.A0(net420),
    .A1(_3933_),
    .S(net85),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _7674_ (.A0(net556),
    .A1(_3934_),
    .S(net85),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _7675_ (.A0(net638),
    .A1(_3935_),
    .S(net85),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _7676_ (.A0(net594),
    .A1(_3936_),
    .S(net85),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _7677_ (.A0(net604),
    .A1(_3937_),
    .S(net85),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _7678_ (.A0(net602),
    .A1(_3938_),
    .S(net85),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _7679_ (.A0(net496),
    .A1(_3939_),
    .S(net85),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _7680_ (.A0(net671),
    .A1(_3940_),
    .S(net85),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _7681_ (.A0(net410),
    .A1(_3941_),
    .S(net85),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _7682_ (.A0(net456),
    .A1(_3942_),
    .S(net85),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _7683_ (.A0(net419),
    .A1(_3943_),
    .S(net86),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _7684_ (.A0(net441),
    .A1(_3944_),
    .S(net85),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _7685_ (.A0(net607),
    .A1(_3945_),
    .S(net86),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _7686_ (.A0(net648),
    .A1(_3946_),
    .S(net86),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _7687_ (.A0(net748),
    .A1(_3947_),
    .S(net86),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _7688_ (.A0(net432),
    .A1(_3948_),
    .S(net86),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _7689_ (.A0(net436),
    .A1(_3949_),
    .S(net86),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _7690_ (.A0(net461),
    .A1(_3950_),
    .S(net86),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _7691_ (.A0(net433),
    .A1(_3951_),
    .S(net85),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _7692_ (.A0(net665),
    .A1(_3952_),
    .S(net85),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _7693_ (.A0(net597),
    .A1(_3953_),
    .S(net85),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _7694_ (.A0(net647),
    .A1(_3954_),
    .S(net85),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _7695_ (.A0(net697),
    .A1(_3955_),
    .S(net85),
    .X(_0196_));
 sky130_fd_sc_hd__a41o_1 _7696_ (.A1(net16),
    .A2(_0561_),
    .A3(net20),
    .A4(_3923_),
    .B1(net31),
    .X(_3957_));
 sky130_fd_sc_hd__mux2_1 _7697_ (.A0(net325),
    .A1(_3925_),
    .S(net84),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _7698_ (.A0(net503),
    .A1(_3926_),
    .S(net84),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _7699_ (.A0(net525),
    .A1(_3927_),
    .S(net84),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _7700_ (.A0(net544),
    .A1(_3928_),
    .S(net84),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _7701_ (.A0(net531),
    .A1(_3929_),
    .S(net84),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _7702_ (.A0(net532),
    .A1(_3930_),
    .S(net84),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _7703_ (.A0(net450),
    .A1(_3931_),
    .S(net84),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _7704_ (.A0(net551),
    .A1(_3932_),
    .S(net84),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _7705_ (.A0(net489),
    .A1(_3933_),
    .S(net83),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _7706_ (.A0(net479),
    .A1(_3934_),
    .S(net83),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _7707_ (.A0(net579),
    .A1(_3935_),
    .S(net83),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _7708_ (.A0(net547),
    .A1(_3936_),
    .S(net83),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _7709_ (.A0(net504),
    .A1(_3937_),
    .S(net83),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _7710_ (.A0(net499),
    .A1(_3938_),
    .S(net83),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _7711_ (.A0(net521),
    .A1(_3939_),
    .S(net83),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _7712_ (.A0(net695),
    .A1(_3940_),
    .S(net83),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _7713_ (.A0(net400),
    .A1(_3941_),
    .S(net83),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _7714_ (.A0(net415),
    .A1(_3942_),
    .S(net83),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _7715_ (.A0(net598),
    .A1(_3943_),
    .S(net84),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _7716_ (.A0(net670),
    .A1(_3944_),
    .S(net83),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _7717_ (.A0(net621),
    .A1(_3945_),
    .S(net84),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _7718_ (.A0(net639),
    .A1(_3946_),
    .S(net84),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _7719_ (.A0(net471),
    .A1(_3947_),
    .S(net84),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _7720_ (.A0(net470),
    .A1(_3948_),
    .S(net84),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _7721_ (.A0(net437),
    .A1(_3949_),
    .S(net84),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _7722_ (.A0(net678),
    .A1(_3950_),
    .S(net84),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _7723_ (.A0(net431),
    .A1(_3951_),
    .S(net83),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _7724_ (.A0(net612),
    .A1(_3952_),
    .S(net83),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _7725_ (.A0(net618),
    .A1(_3953_),
    .S(net83),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _7726_ (.A0(net414),
    .A1(_3954_),
    .S(net83),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _7727_ (.A0(net507),
    .A1(_3955_),
    .S(net83),
    .X(_0227_));
 sky130_fd_sc_hd__a41o_1 _7728_ (.A1(net16),
    .A2(net15),
    .A3(net20),
    .A4(_3923_),
    .B1(net31),
    .X(_3958_));
 sky130_fd_sc_hd__mux2_1 _7729_ (.A0(net341),
    .A1(_3925_),
    .S(net82),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _7730_ (.A0(net445),
    .A1(_3926_),
    .S(net82),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _7731_ (.A0(net500),
    .A1(_3927_),
    .S(net82),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _7732_ (.A0(net502),
    .A1(_3928_),
    .S(net82),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _7733_ (.A0(net512),
    .A1(_3929_),
    .S(net82),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _7734_ (.A0(net535),
    .A1(_3930_),
    .S(net82),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _7735_ (.A0(net476),
    .A1(_3931_),
    .S(net82),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _7736_ (.A0(net523),
    .A1(_3932_),
    .S(net82),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _7737_ (.A0(net407),
    .A1(_3933_),
    .S(net81),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _7738_ (.A0(net582),
    .A1(_3934_),
    .S(net81),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _7739_ (.A0(net605),
    .A1(_3935_),
    .S(net81),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _7740_ (.A0(net567),
    .A1(_3936_),
    .S(net81),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _7741_ (.A0(net472),
    .A1(_3937_),
    .S(net81),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _7742_ (.A0(net546),
    .A1(_3938_),
    .S(net81),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _7743_ (.A0(net528),
    .A1(_3939_),
    .S(net81),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _7744_ (.A0(net667),
    .A1(_3940_),
    .S(net81),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _7745_ (.A0(net515),
    .A1(_3941_),
    .S(net81),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _7746_ (.A0(net495),
    .A1(_3942_),
    .S(net81),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _7747_ (.A0(net491),
    .A1(_3943_),
    .S(net81),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _7748_ (.A0(net728),
    .A1(_3944_),
    .S(net82),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _7749_ (.A0(net590),
    .A1(_3945_),
    .S(net82),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _7750_ (.A0(net600),
    .A1(_3946_),
    .S(net82),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _7751_ (.A0(net465),
    .A1(_3947_),
    .S(net82),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _7752_ (.A0(net427),
    .A1(_3948_),
    .S(net82),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _7753_ (.A0(net413),
    .A1(_3949_),
    .S(net82),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _7754_ (.A0(net454),
    .A1(_3950_),
    .S(net82),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _7755_ (.A0(net626),
    .A1(_3951_),
    .S(net81),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _7756_ (.A0(net707),
    .A1(_3952_),
    .S(net81),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _7757_ (.A0(net645),
    .A1(_3953_),
    .S(net81),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _7758_ (.A0(net448),
    .A1(_3954_),
    .S(net81),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _7759_ (.A0(net389),
    .A1(_3955_),
    .S(net81),
    .X(_0258_));
 sky130_fd_sc_hd__or3b_2 _7760_ (.A(net18),
    .B(_0563_),
    .C_N(net20),
    .X(_3959_));
 sky130_fd_sc_hd__o31ai_1 _7761_ (.A1(net16),
    .A2(net15),
    .A3(_3959_),
    .B1(net210),
    .Y(_3960_));
 sky130_fd_sc_hd__mux2_1 _7762_ (.A0(net387),
    .A1(_3925_),
    .S(net78),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _7763_ (.A0(net494),
    .A1(_3926_),
    .S(net78),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _7764_ (.A0(net536),
    .A1(_3927_),
    .S(net78),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _7765_ (.A0(net565),
    .A1(_3928_),
    .S(net78),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _7766_ (.A0(net541),
    .A1(_3929_),
    .S(net78),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _7767_ (.A0(net552),
    .A1(_3930_),
    .S(net78),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _7768_ (.A0(net444),
    .A1(_3931_),
    .S(net78),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _7769_ (.A0(net572),
    .A1(_3932_),
    .S(net78),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _7770_ (.A0(net423),
    .A1(_3933_),
    .S(net77),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _7771_ (.A0(net591),
    .A1(_3934_),
    .S(net77),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _7772_ (.A0(net596),
    .A1(_3935_),
    .S(net77),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _7773_ (.A0(net585),
    .A1(_3936_),
    .S(net77),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _7774_ (.A0(net558),
    .A1(_3937_),
    .S(net77),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _7775_ (.A0(net571),
    .A1(_3938_),
    .S(net77),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _7776_ (.A0(net616),
    .A1(_3939_),
    .S(net78),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _7777_ (.A0(net684),
    .A1(_3940_),
    .S(net78),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _7778_ (.A0(net412),
    .A1(_3941_),
    .S(net77),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _7779_ (.A0(net439),
    .A1(_3942_),
    .S(net78),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _7780_ (.A0(net603),
    .A1(_3943_),
    .S(net78),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _7781_ (.A0(net691),
    .A1(_3944_),
    .S(net77),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _7782_ (.A0(net589),
    .A1(_3945_),
    .S(net77),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _7783_ (.A0(net451),
    .A1(_3946_),
    .S(net77),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _7784_ (.A0(net468),
    .A1(_3947_),
    .S(net78),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _7785_ (.A0(net485),
    .A1(_3948_),
    .S(net78),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _7786_ (.A0(net438),
    .A1(_3949_),
    .S(net78),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _7787_ (.A0(net622),
    .A1(_3950_),
    .S(net77),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _7788_ (.A0(net474),
    .A1(_3951_),
    .S(net77),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _7789_ (.A0(net628),
    .A1(_3952_),
    .S(net77),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _7790_ (.A0(net674),
    .A1(_3953_),
    .S(net77),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _7791_ (.A0(net505),
    .A1(_3954_),
    .S(net77),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _7792_ (.A0(net623),
    .A1(_3955_),
    .S(net77),
    .X(_0289_));
 sky130_fd_sc_hd__and3_1 _7793_ (.A(_0560_),
    .B(net15),
    .C(net20),
    .X(_3961_));
 sky130_fd_sc_hd__a31o_1 _7794_ (.A1(_0562_),
    .A2(net17),
    .A3(_3961_),
    .B1(net31),
    .X(_3962_));
 sky130_fd_sc_hd__mux2_1 _7795_ (.A0(net347),
    .A1(_3925_),
    .S(net76),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _7796_ (.A0(net526),
    .A1(_3926_),
    .S(net76),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _7797_ (.A0(net518),
    .A1(_3927_),
    .S(net76),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _7798_ (.A0(net570),
    .A1(_3928_),
    .S(net76),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _7799_ (.A0(net524),
    .A1(_3929_),
    .S(net76),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _7800_ (.A0(net562),
    .A1(_3930_),
    .S(net76),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _7801_ (.A0(net466),
    .A1(_3931_),
    .S(net76),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _7802_ (.A0(net555),
    .A1(_3932_),
    .S(net76),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _7803_ (.A0(net430),
    .A1(_3933_),
    .S(net75),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _7804_ (.A0(net553),
    .A1(_3934_),
    .S(net75),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _7805_ (.A0(net563),
    .A1(_3935_),
    .S(net75),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _7806_ (.A0(net569),
    .A1(_3936_),
    .S(net75),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _7807_ (.A0(net506),
    .A1(_3937_),
    .S(net75),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _7808_ (.A0(net595),
    .A1(_3938_),
    .S(net76),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _7809_ (.A0(net601),
    .A1(_3939_),
    .S(net76),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _7810_ (.A0(net681),
    .A1(_3940_),
    .S(net76),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _7811_ (.A0(net440),
    .A1(_3941_),
    .S(net75),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _7812_ (.A0(net527),
    .A1(_3942_),
    .S(net76),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _7813_ (.A0(net615),
    .A1(_3943_),
    .S(net76),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _7814_ (.A0(net629),
    .A1(_3944_),
    .S(net75),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _7815_ (.A0(net539),
    .A1(_3945_),
    .S(net75),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _7816_ (.A0(net557),
    .A1(_3946_),
    .S(net75),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _7817_ (.A0(net422),
    .A1(_3947_),
    .S(net75),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _7818_ (.A0(net480),
    .A1(_3948_),
    .S(net76),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _7819_ (.A0(net447),
    .A1(_3949_),
    .S(net76),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _7820_ (.A0(net701),
    .A1(_3950_),
    .S(net75),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _7821_ (.A0(net534),
    .A1(_3951_),
    .S(net75),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _7822_ (.A0(net624),
    .A1(_3952_),
    .S(net75),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _7823_ (.A0(net609),
    .A1(_3953_),
    .S(net75),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _7824_ (.A0(net404),
    .A1(_3954_),
    .S(net75),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _7825_ (.A0(net559),
    .A1(_3955_),
    .S(net75),
    .X(_0320_));
 sky130_fd_sc_hd__o31ai_1 _7826_ (.A1(_0560_),
    .A2(net15),
    .A3(_3959_),
    .B1(net210),
    .Y(_3963_));
 sky130_fd_sc_hd__mux2_1 _7827_ (.A0(net385),
    .A1(_3925_),
    .S(net74),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _7828_ (.A0(net459),
    .A1(_3926_),
    .S(net74),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _7829_ (.A0(net543),
    .A1(_3927_),
    .S(net74),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _7830_ (.A0(net574),
    .A1(_3928_),
    .S(net74),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _7831_ (.A0(net542),
    .A1(_3929_),
    .S(net74),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _7832_ (.A0(net530),
    .A1(_3930_),
    .S(net74),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _7833_ (.A0(net486),
    .A1(_3931_),
    .S(net74),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _7834_ (.A0(net578),
    .A1(_3932_),
    .S(net74),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _7835_ (.A0(net337),
    .A1(_3933_),
    .S(net73),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _7836_ (.A0(net488),
    .A1(_3934_),
    .S(net73),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _7837_ (.A0(net421),
    .A1(_3935_),
    .S(net73),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _7838_ (.A0(net484),
    .A1(_3936_),
    .S(net73),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _7839_ (.A0(net408),
    .A1(_3937_),
    .S(net73),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _7840_ (.A0(net614),
    .A1(_3938_),
    .S(net73),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _7841_ (.A0(net588),
    .A1(_3939_),
    .S(net74),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _7842_ (.A0(net677),
    .A1(_3940_),
    .S(net74),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _7843_ (.A0(net369),
    .A1(_3941_),
    .S(net73),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _7844_ (.A0(net335),
    .A1(_3942_),
    .S(net73),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _7845_ (.A0(net463),
    .A1(_3943_),
    .S(net73),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _7846_ (.A0(net655),
    .A1(_3944_),
    .S(net73),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _7847_ (.A0(net651),
    .A1(_3945_),
    .S(net73),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _7848_ (.A0(net475),
    .A1(_3946_),
    .S(net73),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _7849_ (.A0(net399),
    .A1(_3947_),
    .S(net73),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _7850_ (.A0(net493),
    .A1(_3948_),
    .S(net74),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _7851_ (.A0(net446),
    .A1(_3949_),
    .S(net74),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _7852_ (.A0(net529),
    .A1(_3950_),
    .S(net74),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _7853_ (.A0(net487),
    .A1(_3951_),
    .S(net74),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _7854_ (.A0(net481),
    .A1(_3952_),
    .S(net74),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _7855_ (.A0(net568),
    .A1(_3953_),
    .S(net73),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _7856_ (.A0(net498),
    .A1(_3954_),
    .S(net73),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _7857_ (.A0(net321),
    .A1(_3955_),
    .S(net73),
    .X(_0351_));
 sky130_fd_sc_hd__o31ai_2 _7858_ (.A1(_0560_),
    .A2(_0561_),
    .A3(_3959_),
    .B1(net210),
    .Y(_3964_));
 sky130_fd_sc_hd__mux2_1 _7859_ (.A0(net367),
    .A1(_3925_),
    .S(net72),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _7860_ (.A0(net511),
    .A1(_3926_),
    .S(net72),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _7861_ (.A0(net514),
    .A1(_3927_),
    .S(net72),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _7862_ (.A0(net554),
    .A1(_3928_),
    .S(net72),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _7863_ (.A0(net516),
    .A1(_3929_),
    .S(net72),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _7864_ (.A0(net509),
    .A1(_3930_),
    .S(net72),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _7865_ (.A0(net460),
    .A1(_3931_),
    .S(net72),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _7866_ (.A0(net564),
    .A1(_3932_),
    .S(net72),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _7867_ (.A0(net497),
    .A1(_3933_),
    .S(net71),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _7868_ (.A0(net469),
    .A1(_3934_),
    .S(net71),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _7869_ (.A0(net508),
    .A1(_3935_),
    .S(net71),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _7870_ (.A0(net458),
    .A1(_3936_),
    .S(net71),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _7871_ (.A0(net443),
    .A1(_3937_),
    .S(net71),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _7872_ (.A0(net575),
    .A1(_3938_),
    .S(net71),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _7873_ (.A0(net592),
    .A1(_3939_),
    .S(net72),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _7874_ (.A0(net687),
    .A1(_3940_),
    .S(net72),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _7875_ (.A0(net538),
    .A1(_3941_),
    .S(net71),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _7876_ (.A0(net637),
    .A1(_3942_),
    .S(net72),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _7877_ (.A0(net679),
    .A1(_3943_),
    .S(net72),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _7878_ (.A0(net641),
    .A1(_3944_),
    .S(net71),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _7879_ (.A0(net663),
    .A1(_3945_),
    .S(net71),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _7880_ (.A0(net633),
    .A1(_3946_),
    .S(net71),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _7881_ (.A0(net483),
    .A1(_3947_),
    .S(net71),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _7882_ (.A0(net424),
    .A1(_3948_),
    .S(net72),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _7883_ (.A0(net428),
    .A1(_3949_),
    .S(net72),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _7884_ (.A0(net425),
    .A1(_3950_),
    .S(net72),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _7885_ (.A0(net501),
    .A1(_3951_),
    .S(net71),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _7886_ (.A0(net627),
    .A1(_3952_),
    .S(net71),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _7887_ (.A0(net593),
    .A1(_3953_),
    .S(net71),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _7888_ (.A0(net640),
    .A1(_3954_),
    .S(net71),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _7889_ (.A0(net613),
    .A1(_3955_),
    .S(net71),
    .X(_0382_));
 sky130_fd_sc_hd__nor2_1 _7890_ (.A(net16),
    .B(net15),
    .Y(_3965_));
 sky130_fd_sc_hd__a41o_1 _7891_ (.A1(net18),
    .A2(_0563_),
    .A3(net20),
    .A4(_3965_),
    .B1(net31),
    .X(_3966_));
 sky130_fd_sc_hd__mux2_1 _7892_ (.A0(net381),
    .A1(_3925_),
    .S(net80),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _7893_ (.A0(net417),
    .A1(_3926_),
    .S(net80),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _7894_ (.A0(net513),
    .A1(_3927_),
    .S(net80),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _7895_ (.A0(net560),
    .A1(_3928_),
    .S(net80),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _7896_ (.A0(net492),
    .A1(_3929_),
    .S(net80),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _7897_ (.A0(net550),
    .A1(_3930_),
    .S(net80),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _7898_ (.A0(net580),
    .A1(_3931_),
    .S(net80),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _7899_ (.A0(net533),
    .A1(_3932_),
    .S(net80),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _7900_ (.A0(net545),
    .A1(_3933_),
    .S(net79),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _7901_ (.A0(net426),
    .A1(_3934_),
    .S(net79),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _7902_ (.A0(net442),
    .A1(_3935_),
    .S(net79),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _7903_ (.A0(net435),
    .A1(_3936_),
    .S(net79),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _7904_ (.A0(net490),
    .A1(_3937_),
    .S(net79),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _7905_ (.A0(net519),
    .A1(_3938_),
    .S(net79),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _7906_ (.A0(net583),
    .A1(_3939_),
    .S(net79),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _7907_ (.A0(net669),
    .A1(_3940_),
    .S(net79),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _7908_ (.A0(net464),
    .A1(_3941_),
    .S(net79),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _7909_ (.A0(net587),
    .A1(_3942_),
    .S(net79),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _7910_ (.A0(net708),
    .A1(_3943_),
    .S(net80),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _7911_ (.A0(net646),
    .A1(_3944_),
    .S(net79),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _7912_ (.A0(net634),
    .A1(_3945_),
    .S(net79),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _7913_ (.A0(net632),
    .A1(_3946_),
    .S(net79),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _7914_ (.A0(net478),
    .A1(_3947_),
    .S(net80),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _7915_ (.A0(net418),
    .A1(_3948_),
    .S(net80),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _7916_ (.A0(net411),
    .A1(_3949_),
    .S(net80),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _7917_ (.A0(net517),
    .A1(_3950_),
    .S(net80),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _7918_ (.A0(net455),
    .A1(_3951_),
    .S(net80),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _7919_ (.A0(net643),
    .A1(_3952_),
    .S(net80),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _7920_ (.A0(net586),
    .A1(_3953_),
    .S(net79),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _7921_ (.A0(net676),
    .A1(_3954_),
    .S(net79),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _7922_ (.A0(net610),
    .A1(_3955_),
    .S(net79),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _7923_ (.A0(net718),
    .A1(\ann.sum[0] ),
    .S(net65),
    .X(_3967_));
 sky130_fd_sc_hd__and2_1 _7924_ (.A(net201),
    .B(_3967_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _7925_ (.A0(net736),
    .A1(\ann.sum[1] ),
    .S(net65),
    .X(_3968_));
 sky130_fd_sc_hd__and2_1 _7926_ (.A(net201),
    .B(_3968_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _7927_ (.A0(net737),
    .A1(\ann.sum[2] ),
    .S(net64),
    .X(_3969_));
 sky130_fd_sc_hd__and2_1 _7928_ (.A(net201),
    .B(_3969_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _7929_ (.A0(net729),
    .A1(\ann.sum[3] ),
    .S(net65),
    .X(_3970_));
 sky130_fd_sc_hd__and2_1 _7930_ (.A(net204),
    .B(_3970_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _7931_ (.A0(net720),
    .A1(\ann.sum[4] ),
    .S(net64),
    .X(_3971_));
 sky130_fd_sc_hd__and2_1 _7932_ (.A(net203),
    .B(_3971_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _7933_ (.A0(net781),
    .A1(\ann.sum[5] ),
    .S(net64),
    .X(_3972_));
 sky130_fd_sc_hd__and2_1 _7934_ (.A(net204),
    .B(_3972_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _7935_ (.A0(net763),
    .A1(\ann.sum[6] ),
    .S(net64),
    .X(_3973_));
 sky130_fd_sc_hd__and2_1 _7936_ (.A(net203),
    .B(_3973_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _7937_ (.A0(net739),
    .A1(\ann.sum[7] ),
    .S(net65),
    .X(_3974_));
 sky130_fd_sc_hd__and2_1 _7938_ (.A(net203),
    .B(_3974_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _7939_ (.A0(net733),
    .A1(\ann.sum[8] ),
    .S(net65),
    .X(_3975_));
 sky130_fd_sc_hd__and2_1 _7940_ (.A(net206),
    .B(_3975_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _7941_ (.A0(net723),
    .A1(\ann.sum[9] ),
    .S(net65),
    .X(_3976_));
 sky130_fd_sc_hd__and2_1 _7942_ (.A(net205),
    .B(_3976_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _7943_ (.A0(net715),
    .A1(\ann.sum[10] ),
    .S(net65),
    .X(_3977_));
 sky130_fd_sc_hd__and2_1 _7944_ (.A(net205),
    .B(_3977_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _7945_ (.A0(net767),
    .A1(\ann.sum[11] ),
    .S(net65),
    .X(_3978_));
 sky130_fd_sc_hd__and2_1 _7946_ (.A(net205),
    .B(_3978_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _7947_ (.A0(net752),
    .A1(\ann.sum[12] ),
    .S(net65),
    .X(_3979_));
 sky130_fd_sc_hd__and2_1 _7948_ (.A(net205),
    .B(_3979_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _7949_ (.A0(net766),
    .A1(\ann.sum[13] ),
    .S(net65),
    .X(_3980_));
 sky130_fd_sc_hd__and2_1 _7950_ (.A(net207),
    .B(_3980_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _7951_ (.A0(net746),
    .A1(\ann.sum[14] ),
    .S(net65),
    .X(_3981_));
 sky130_fd_sc_hd__and2_1 _7952_ (.A(net202),
    .B(_3981_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _7953_ (.A0(net719),
    .A1(\ann.sum[15] ),
    .S(net65),
    .X(_3982_));
 sky130_fd_sc_hd__and2_1 _7954_ (.A(net202),
    .B(_3982_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _7955_ (.A0(net741),
    .A1(\ann.sum[16] ),
    .S(net65),
    .X(_3983_));
 sky130_fd_sc_hd__and2_1 _7956_ (.A(net201),
    .B(_3983_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _7957_ (.A0(net721),
    .A1(\ann.sum[17] ),
    .S(net64),
    .X(_3984_));
 sky130_fd_sc_hd__and2_1 _7958_ (.A(net201),
    .B(_3984_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _7959_ (.A0(net714),
    .A1(\ann.sum[18] ),
    .S(net65),
    .X(_3985_));
 sky130_fd_sc_hd__and2_1 _7960_ (.A(net199),
    .B(_3985_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _7961_ (.A0(net738),
    .A1(\ann.sum[19] ),
    .S(net64),
    .X(_3986_));
 sky130_fd_sc_hd__and2_1 _7962_ (.A(net199),
    .B(_3986_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _7963_ (.A0(net768),
    .A1(\ann.sum[20] ),
    .S(net64),
    .X(_3987_));
 sky130_fd_sc_hd__and2_1 _7964_ (.A(net197),
    .B(_3987_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _7965_ (.A0(net777),
    .A1(\ann.sum[21] ),
    .S(net64),
    .X(_3988_));
 sky130_fd_sc_hd__and2_1 _7966_ (.A(net197),
    .B(_3988_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _7967_ (.A0(net751),
    .A1(\ann.sum[22] ),
    .S(net64),
    .X(_3989_));
 sky130_fd_sc_hd__and2_1 _7968_ (.A(net200),
    .B(_3989_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _7969_ (.A0(net726),
    .A1(\ann.sum[23] ),
    .S(net64),
    .X(_3990_));
 sky130_fd_sc_hd__and2_1 _7970_ (.A(net197),
    .B(_3990_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _7971_ (.A0(net769),
    .A1(\ann.sum[24] ),
    .S(net64),
    .X(_3991_));
 sky130_fd_sc_hd__and2_1 _7972_ (.A(net196),
    .B(_3991_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _7973_ (.A0(net776),
    .A1(\ann.sum[25] ),
    .S(net64),
    .X(_3992_));
 sky130_fd_sc_hd__and2_1 _7974_ (.A(net196),
    .B(_3992_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _7975_ (.A0(net722),
    .A1(\ann.sum[26] ),
    .S(net64),
    .X(_3993_));
 sky130_fd_sc_hd__and2_1 _7976_ (.A(net196),
    .B(_3993_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _7977_ (.A0(net756),
    .A1(\ann.sum[27] ),
    .S(net64),
    .X(_3994_));
 sky130_fd_sc_hd__and2_1 _7978_ (.A(net196),
    .B(_3994_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _7979_ (.A0(net705),
    .A1(\ann.sum[28] ),
    .S(net64),
    .X(_3995_));
 sky130_fd_sc_hd__and2_1 _7980_ (.A(net198),
    .B(_3995_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _7981_ (.A0(net713),
    .A1(\ann.sum[29] ),
    .S(net64),
    .X(_3996_));
 sky130_fd_sc_hd__and2_1 _7982_ (.A(net198),
    .B(_3996_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _7983_ (.A0(net716),
    .A1(\ann.sum[30] ),
    .S(\ann.ldX ),
    .X(_3997_));
 sky130_fd_sc_hd__and2_1 _7984_ (.A(net199),
    .B(_3997_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _7985_ (.A0(net702),
    .A1(net59),
    .S(net65),
    .X(_3998_));
 sky130_fd_sc_hd__and2_1 _7986_ (.A(net198),
    .B(_3998_),
    .X(_0445_));
 sky130_fd_sc_hd__a31o_1 _7987_ (.A1(net18),
    .A2(_0563_),
    .A3(_3961_),
    .B1(net31),
    .X(_3999_));
 sky130_fd_sc_hd__mux2_1 _7988_ (.A0(net393),
    .A1(_3925_),
    .S(net70),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _7989_ (.A0(net449),
    .A1(_3926_),
    .S(net70),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _7990_ (.A0(net577),
    .A1(_3927_),
    .S(net70),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _7991_ (.A0(net482),
    .A1(_3928_),
    .S(net70),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _7992_ (.A0(net606),
    .A1(_3929_),
    .S(net70),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _7993_ (.A0(net549),
    .A1(_3930_),
    .S(net70),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _7994_ (.A0(net477),
    .A1(_3931_),
    .S(net70),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _7995_ (.A0(net576),
    .A1(_3932_),
    .S(net70),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _7996_ (.A0(net429),
    .A1(_3933_),
    .S(net69),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _7997_ (.A0(net434),
    .A1(_3934_),
    .S(net69),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _7998_ (.A0(net510),
    .A1(_3935_),
    .S(net69),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _7999_ (.A0(net473),
    .A1(_3936_),
    .S(net69),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _8000_ (.A0(net620),
    .A1(_3937_),
    .S(net69),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _8001_ (.A0(net650),
    .A1(_3938_),
    .S(net69),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _8002_ (.A0(net617),
    .A1(_3939_),
    .S(net69),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _8003_ (.A0(net682),
    .A1(_3940_),
    .S(net69),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _8004_ (.A0(net452),
    .A1(_3941_),
    .S(net69),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _8005_ (.A0(net406),
    .A1(_3942_),
    .S(net69),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _8006_ (.A0(net636),
    .A1(_3943_),
    .S(net69),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _8007_ (.A0(net673),
    .A1(_3944_),
    .S(net69),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _8008_ (.A0(net659),
    .A1(_3945_),
    .S(net69),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _8009_ (.A0(net599),
    .A1(_3946_),
    .S(net70),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _8010_ (.A0(net657),
    .A1(_3947_),
    .S(net70),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _8011_ (.A0(net453),
    .A1(_3948_),
    .S(net70),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _8012_ (.A0(net548),
    .A1(_3949_),
    .S(net70),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _8013_ (.A0(net608),
    .A1(_3950_),
    .S(net70),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _8014_ (.A0(net581),
    .A1(_3951_),
    .S(net70),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _8015_ (.A0(net664),
    .A1(_3952_),
    .S(net70),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _8016_ (.A0(net462),
    .A1(_3953_),
    .S(net69),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _8017_ (.A0(net672),
    .A1(_3954_),
    .S(net69),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _8018_ (.A0(net631),
    .A1(_3955_),
    .S(net69),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _8019_ (.A0(net783),
    .A1(net29),
    .S(net22),
    .X(_4000_));
 sky130_fd_sc_hd__and2_1 _8020_ (.A(net210),
    .B(_4000_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _8021_ (.A0(net754),
    .A1(net30),
    .S(net22),
    .X(_4001_));
 sky130_fd_sc_hd__and2_1 _8022_ (.A(net210),
    .B(_4001_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _8023_ (.A0(net704),
    .A1(net1),
    .S(net22),
    .X(_4002_));
 sky130_fd_sc_hd__and2_1 _8024_ (.A(net215),
    .B(_4002_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _8025_ (.A0(net724),
    .A1(net2),
    .S(net22),
    .X(_4003_));
 sky130_fd_sc_hd__and2_1 _8026_ (.A(net215),
    .B(_4003_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _8027_ (.A0(net734),
    .A1(net3),
    .S(net22),
    .X(_4004_));
 sky130_fd_sc_hd__and2_1 _8028_ (.A(net210),
    .B(_4004_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _8029_ (.A0(net711),
    .A1(net4),
    .S(net22),
    .X(_4005_));
 sky130_fd_sc_hd__and2_1 _8030_ (.A(net215),
    .B(_4005_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _8031_ (.A0(net770),
    .A1(net5),
    .S(net22),
    .X(_4006_));
 sky130_fd_sc_hd__and2_1 _8032_ (.A(net215),
    .B(_4006_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _8033_ (.A0(net762),
    .A1(net6),
    .S(net22),
    .X(_4007_));
 sky130_fd_sc_hd__and2_1 _8034_ (.A(net215),
    .B(_4007_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _8035_ (.A0(net779),
    .A1(net7),
    .S(net22),
    .X(_4008_));
 sky130_fd_sc_hd__and2_1 _8036_ (.A(net215),
    .B(_4008_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _8037_ (.A0(net775),
    .A1(net8),
    .S(net22),
    .X(_4009_));
 sky130_fd_sc_hd__and2_1 _8038_ (.A(net215),
    .B(_4009_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _8039_ (.A0(net786),
    .A1(net9),
    .S(net22),
    .X(_4010_));
 sky130_fd_sc_hd__and2_1 _8040_ (.A(net210),
    .B(_4010_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _8041_ (.A0(net787),
    .A1(net10),
    .S(net22),
    .X(_4011_));
 sky130_fd_sc_hd__and2_1 _8042_ (.A(net211),
    .B(_4011_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _8043_ (.A0(net740),
    .A1(net11),
    .S(net22),
    .X(_4012_));
 sky130_fd_sc_hd__and2_1 _8044_ (.A(net210),
    .B(_4012_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _8045_ (.A0(net780),
    .A1(net12),
    .S(net22),
    .X(_4013_));
 sky130_fd_sc_hd__and2_1 _8046_ (.A(net211),
    .B(_4013_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _8047_ (.A0(net742),
    .A1(net13),
    .S(net22),
    .X(_4014_));
 sky130_fd_sc_hd__and2_1 _8048_ (.A(net211),
    .B(_4014_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _8049_ (.A0(net735),
    .A1(net14),
    .S(net22),
    .X(_4015_));
 sky130_fd_sc_hd__and2_1 _8050_ (.A(net211),
    .B(_4015_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _8051_ (.A0(net778),
    .A1(net29),
    .S(net23),
    .X(_4016_));
 sky130_fd_sc_hd__and2_1 _8052_ (.A(net210),
    .B(_4016_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _8053_ (.A0(net745),
    .A1(net30),
    .S(net23),
    .X(_4017_));
 sky130_fd_sc_hd__and2_1 _8054_ (.A(net210),
    .B(_4017_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _8055_ (.A0(net759),
    .A1(net1),
    .S(net23),
    .X(_4018_));
 sky130_fd_sc_hd__and2_1 _8056_ (.A(net210),
    .B(_4018_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _8057_ (.A0(net725),
    .A1(net2),
    .S(net23),
    .X(_4019_));
 sky130_fd_sc_hd__and2_1 _8058_ (.A(net210),
    .B(_4019_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _8059_ (.A0(net761),
    .A1(net3),
    .S(net23),
    .X(_4020_));
 sky130_fd_sc_hd__and2_1 _8060_ (.A(net210),
    .B(_4020_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _8061_ (.A0(net764),
    .A1(net4),
    .S(net23),
    .X(_4021_));
 sky130_fd_sc_hd__and2_1 _8062_ (.A(net210),
    .B(_4021_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _8063_ (.A0(net710),
    .A1(net5),
    .S(net23),
    .X(_4022_));
 sky130_fd_sc_hd__and2_1 _8064_ (.A(net210),
    .B(_4022_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _8065_ (.A0(net730),
    .A1(net6),
    .S(net23),
    .X(_4023_));
 sky130_fd_sc_hd__and2_1 _8066_ (.A(net215),
    .B(_4023_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _8067_ (.A0(net760),
    .A1(net7),
    .S(net23),
    .X(_4024_));
 sky130_fd_sc_hd__and2_1 _8068_ (.A(net212),
    .B(_4024_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _8069_ (.A0(net709),
    .A1(net8),
    .S(net23),
    .X(_4025_));
 sky130_fd_sc_hd__and2_1 _8070_ (.A(net212),
    .B(_4025_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _8071_ (.A0(net744),
    .A1(net9),
    .S(net23),
    .X(_4026_));
 sky130_fd_sc_hd__and2_1 _8072_ (.A(net212),
    .B(_4026_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _8073_ (.A0(net732),
    .A1(net10),
    .S(net23),
    .X(_4027_));
 sky130_fd_sc_hd__and2_1 _8074_ (.A(net212),
    .B(_4027_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _8075_ (.A0(net727),
    .A1(net11),
    .S(net23),
    .X(_4028_));
 sky130_fd_sc_hd__and2_1 _8076_ (.A(net212),
    .B(_4028_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _8077_ (.A0(net771),
    .A1(net12),
    .S(net23),
    .X(_4029_));
 sky130_fd_sc_hd__and2_1 _8078_ (.A(net211),
    .B(_4029_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _8079_ (.A0(net772),
    .A1(net13),
    .S(net23),
    .X(_4030_));
 sky130_fd_sc_hd__and2_1 _8080_ (.A(net211),
    .B(_4030_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _8081_ (.A0(net749),
    .A1(net14),
    .S(net23),
    .X(_4031_));
 sky130_fd_sc_hd__and2_1 _8082_ (.A(net211),
    .B(_4031_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _8083_ (.A0(net680),
    .A1(net145),
    .S(net218),
    .X(_4032_));
 sky130_fd_sc_hd__nand2b_1 _8084_ (.A_N(net29),
    .B(net216),
    .Y(_4033_));
 sky130_fd_sc_hd__o211a_1 _8085_ (.A1(net216),
    .A2(_4032_),
    .B1(_4033_),
    .C1(net211),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _8086_ (.A0(net683),
    .A1(net143),
    .S(net218),
    .X(_4034_));
 sky130_fd_sc_hd__nand2b_1 _8087_ (.A_N(net30),
    .B(net216),
    .Y(_4035_));
 sky130_fd_sc_hd__o211a_1 _8088_ (.A1(net216),
    .A2(_4034_),
    .B1(_4035_),
    .C1(net211),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _8089_ (.A0(net688),
    .A1(net140),
    .S(net218),
    .X(_4036_));
 sky130_fd_sc_hd__nand2b_1 _8090_ (.A_N(net1),
    .B(net216),
    .Y(_4037_));
 sky130_fd_sc_hd__o211a_1 _8091_ (.A1(net216),
    .A2(_4036_),
    .B1(_4037_),
    .C1(net211),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _8092_ (.A0(net686),
    .A1(net137),
    .S(net218),
    .X(_4038_));
 sky130_fd_sc_hd__nand2b_1 _8093_ (.A_N(net2),
    .B(net216),
    .Y(_4039_));
 sky130_fd_sc_hd__o211a_1 _8094_ (.A1(net216),
    .A2(_4038_),
    .B1(_4039_),
    .C1(net211),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _8095_ (.A0(net692),
    .A1(net134),
    .S(net218),
    .X(_4040_));
 sky130_fd_sc_hd__nand2b_1 _8096_ (.A_N(net3),
    .B(net217),
    .Y(_4041_));
 sky130_fd_sc_hd__o211a_1 _8097_ (.A1(net217),
    .A2(_4040_),
    .B1(_4041_),
    .C1(net213),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _8098_ (.A0(net694),
    .A1(net131),
    .S(net218),
    .X(_4042_));
 sky130_fd_sc_hd__nand2b_1 _8099_ (.A_N(net4),
    .B(net217),
    .Y(_4043_));
 sky130_fd_sc_hd__o211a_1 _8100_ (.A1(net217),
    .A2(_4042_),
    .B1(_4043_),
    .C1(net213),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _8101_ (.A0(net690),
    .A1(net128),
    .S(net218),
    .X(_4044_));
 sky130_fd_sc_hd__nand2b_1 _8102_ (.A_N(net5),
    .B(net217),
    .Y(_4045_));
 sky130_fd_sc_hd__o211a_1 _8103_ (.A1(net217),
    .A2(_4044_),
    .B1(_4045_),
    .C1(net213),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _8104_ (.A0(net689),
    .A1(net126),
    .S(net218),
    .X(_4046_));
 sky130_fd_sc_hd__nand2b_1 _8105_ (.A_N(net6),
    .B(net217),
    .Y(_4047_));
 sky130_fd_sc_hd__o211a_1 _8106_ (.A1(net217),
    .A2(_4046_),
    .B1(_4047_),
    .C1(net213),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _8107_ (.A0(net693),
    .A1(net124),
    .S(net218),
    .X(_4048_));
 sky130_fd_sc_hd__nand2b_1 _8108_ (.A_N(net7),
    .B(net217),
    .Y(_4049_));
 sky130_fd_sc_hd__o211a_1 _8109_ (.A1(net217),
    .A2(_4048_),
    .B1(_4049_),
    .C1(net214),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _8110_ (.A0(net685),
    .A1(net122),
    .S(net218),
    .X(_4050_));
 sky130_fd_sc_hd__nand2b_1 _8111_ (.A_N(net8),
    .B(net217),
    .Y(_4051_));
 sky130_fd_sc_hd__o211a_1 _8112_ (.A1(net217),
    .A2(_4050_),
    .B1(_4051_),
    .C1(net213),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _8113_ (.A0(net699),
    .A1(net119),
    .S(net218),
    .X(_4052_));
 sky130_fd_sc_hd__nand2b_1 _8114_ (.A_N(net9),
    .B(net217),
    .Y(_4053_));
 sky130_fd_sc_hd__o211a_1 _8115_ (.A1(net27),
    .A2(_4052_),
    .B1(_4053_),
    .C1(net213),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _8116_ (.A0(net698),
    .A1(net116),
    .S(net218),
    .X(_4054_));
 sky130_fd_sc_hd__nand2b_1 _8117_ (.A_N(net10),
    .B(net216),
    .Y(_4055_));
 sky130_fd_sc_hd__o211a_1 _8118_ (.A1(net216),
    .A2(_4054_),
    .B1(_4055_),
    .C1(net211),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _8119_ (.A0(net700),
    .A1(net113),
    .S(net25),
    .X(_4056_));
 sky130_fd_sc_hd__nand2b_1 _8120_ (.A_N(net11),
    .B(net27),
    .Y(_4057_));
 sky130_fd_sc_hd__o211a_1 _8121_ (.A1(net27),
    .A2(_4056_),
    .B1(_4057_),
    .C1(net213),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _8122_ (.A0(net706),
    .A1(net110),
    .S(net218),
    .X(_4058_));
 sky130_fd_sc_hd__nand2b_1 _8123_ (.A_N(net12),
    .B(net216),
    .Y(_4059_));
 sky130_fd_sc_hd__o211a_1 _8124_ (.A1(net216),
    .A2(_4058_),
    .B1(_4059_),
    .C1(net211),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _8125_ (.A0(net696),
    .A1(net108),
    .S(net218),
    .X(_4060_));
 sky130_fd_sc_hd__nand2b_1 _8126_ (.A_N(net13),
    .B(net216),
    .Y(_4061_));
 sky130_fd_sc_hd__o211a_1 _8127_ (.A1(net216),
    .A2(_4060_),
    .B1(_4061_),
    .C1(net212),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _8128_ (.A0(net703),
    .A1(net106),
    .S(net25),
    .X(_4062_));
 sky130_fd_sc_hd__nand2b_1 _8129_ (.A_N(net14),
    .B(net217),
    .Y(_4063_));
 sky130_fd_sc_hd__o211a_1 _8130_ (.A1(net217),
    .A2(_4062_),
    .B1(_4063_),
    .C1(net213),
    .X(_0524_));
 sky130_fd_sc_hd__nor2_1 _8131_ (.A(net216),
    .B(net218),
    .Y(_4064_));
 sky130_fd_sc_hd__or2_1 _8132_ (.A(net216),
    .B(net218),
    .X(_4065_));
 sky130_fd_sc_hd__or2_1 _8133_ (.A(\ann.in_ff[0][0] ),
    .B(net192),
    .X(_4066_));
 sky130_fd_sc_hd__o211a_1 _8134_ (.A1(net331),
    .A2(net190),
    .B1(_4066_),
    .C1(net212),
    .X(_0525_));
 sky130_fd_sc_hd__or2_1 _8135_ (.A(\ann.in_ff[0][1] ),
    .B(net192),
    .X(_4067_));
 sky130_fd_sc_hd__o211a_1 _8136_ (.A1(net345),
    .A2(net190),
    .B1(_4067_),
    .C1(net212),
    .X(_0526_));
 sky130_fd_sc_hd__or2_1 _8137_ (.A(net688),
    .B(net192),
    .X(_4068_));
 sky130_fd_sc_hd__o211a_1 _8138_ (.A1(net371),
    .A2(net190),
    .B1(_4068_),
    .C1(net212),
    .X(_0527_));
 sky130_fd_sc_hd__or2_1 _8139_ (.A(net686),
    .B(net192),
    .X(_4069_));
 sky130_fd_sc_hd__o211a_1 _8140_ (.A1(net373),
    .A2(net190),
    .B1(_4069_),
    .C1(net213),
    .X(_0528_));
 sky130_fd_sc_hd__or2_1 _8141_ (.A(\ann.in_ff[0][4] ),
    .B(net193),
    .X(_4070_));
 sky130_fd_sc_hd__o211a_1 _8142_ (.A1(net361),
    .A2(net191),
    .B1(_4070_),
    .C1(net214),
    .X(_0529_));
 sky130_fd_sc_hd__or2_1 _8143_ (.A(\ann.in_ff[0][5] ),
    .B(net193),
    .X(_4071_));
 sky130_fd_sc_hd__o211a_1 _8144_ (.A1(net363),
    .A2(net191),
    .B1(_4071_),
    .C1(net214),
    .X(_0530_));
 sky130_fd_sc_hd__or2_1 _8145_ (.A(\ann.in_ff[0][6] ),
    .B(net193),
    .X(_4072_));
 sky130_fd_sc_hd__o211a_1 _8146_ (.A1(net375),
    .A2(net191),
    .B1(_4072_),
    .C1(net214),
    .X(_0531_));
 sky130_fd_sc_hd__or2_1 _8147_ (.A(net689),
    .B(net193),
    .X(_4073_));
 sky130_fd_sc_hd__o211a_1 _8148_ (.A1(net327),
    .A2(net191),
    .B1(_4073_),
    .C1(net214),
    .X(_0532_));
 sky130_fd_sc_hd__or2_1 _8149_ (.A(\ann.in_ff[0][8] ),
    .B(net193),
    .X(_4074_));
 sky130_fd_sc_hd__o211a_1 _8150_ (.A1(net359),
    .A2(net191),
    .B1(_4074_),
    .C1(net214),
    .X(_0533_));
 sky130_fd_sc_hd__or2_1 _8151_ (.A(\ann.in_ff[0][9] ),
    .B(net193),
    .X(_4075_));
 sky130_fd_sc_hd__o211a_1 _8152_ (.A1(net377),
    .A2(net191),
    .B1(_4075_),
    .C1(net214),
    .X(_0534_));
 sky130_fd_sc_hd__or2_1 _8153_ (.A(\ann.in_ff[0][10] ),
    .B(net193),
    .X(_4076_));
 sky130_fd_sc_hd__o211a_1 _8154_ (.A1(net391),
    .A2(net191),
    .B1(_4076_),
    .C1(net213),
    .X(_0535_));
 sky130_fd_sc_hd__or2_1 _8155_ (.A(\ann.in_ff[0][11] ),
    .B(net192),
    .X(_4077_));
 sky130_fd_sc_hd__o211a_1 _8156_ (.A1(net395),
    .A2(net190),
    .B1(_4077_),
    .C1(net212),
    .X(_0536_));
 sky130_fd_sc_hd__or2_1 _8157_ (.A(\ann.in_ff[0][12] ),
    .B(net193),
    .X(_4078_));
 sky130_fd_sc_hd__o211a_1 _8158_ (.A1(net357),
    .A2(net191),
    .B1(_4078_),
    .C1(net213),
    .X(_0537_));
 sky130_fd_sc_hd__or2_1 _8159_ (.A(\ann.in_ff[0][13] ),
    .B(net192),
    .X(_4079_));
 sky130_fd_sc_hd__o211a_1 _8160_ (.A1(net397),
    .A2(net190),
    .B1(_4079_),
    .C1(net211),
    .X(_0538_));
 sky130_fd_sc_hd__or2_1 _8161_ (.A(\ann.in_ff[0][14] ),
    .B(net192),
    .X(_4080_));
 sky130_fd_sc_hd__o211a_1 _8162_ (.A1(net355),
    .A2(net190),
    .B1(_4080_),
    .C1(net211),
    .X(_0539_));
 sky130_fd_sc_hd__or2_1 _8163_ (.A(\ann.in_ff[0][15] ),
    .B(net192),
    .X(_4081_));
 sky130_fd_sc_hd__o211a_1 _8164_ (.A1(net383),
    .A2(net190),
    .B1(_4081_),
    .C1(net213),
    .X(_0540_));
 sky130_fd_sc_hd__or2_1 _8165_ (.A(net331),
    .B(net192),
    .X(_4082_));
 sky130_fd_sc_hd__o211a_1 _8166_ (.A1(net145),
    .A2(net190),
    .B1(_4082_),
    .C1(net212),
    .X(_0541_));
 sky130_fd_sc_hd__or2_1 _8167_ (.A(net345),
    .B(net192),
    .X(_4083_));
 sky130_fd_sc_hd__o211a_1 _8168_ (.A1(net143),
    .A2(net190),
    .B1(_4083_),
    .C1(net212),
    .X(_0542_));
 sky130_fd_sc_hd__or2_1 _8169_ (.A(net371),
    .B(net192),
    .X(_4084_));
 sky130_fd_sc_hd__o211a_1 _8170_ (.A1(net140),
    .A2(net190),
    .B1(_4084_),
    .C1(net212),
    .X(_0543_));
 sky130_fd_sc_hd__or2_1 _8171_ (.A(net373),
    .B(net192),
    .X(_4085_));
 sky130_fd_sc_hd__o211a_1 _8172_ (.A1(net137),
    .A2(net190),
    .B1(_4085_),
    .C1(net214),
    .X(_0544_));
 sky130_fd_sc_hd__or2_1 _8173_ (.A(net361),
    .B(net193),
    .X(_4086_));
 sky130_fd_sc_hd__o211a_1 _8174_ (.A1(net134),
    .A2(net191),
    .B1(_4086_),
    .C1(net214),
    .X(_0545_));
 sky130_fd_sc_hd__or2_1 _8175_ (.A(net363),
    .B(net193),
    .X(_4087_));
 sky130_fd_sc_hd__o211a_1 _8176_ (.A1(net131),
    .A2(net191),
    .B1(_4087_),
    .C1(net214),
    .X(_0546_));
 sky130_fd_sc_hd__or2_1 _8177_ (.A(net375),
    .B(net193),
    .X(_4088_));
 sky130_fd_sc_hd__o211a_1 _8178_ (.A1(net128),
    .A2(net191),
    .B1(_4088_),
    .C1(net214),
    .X(_0547_));
 sky130_fd_sc_hd__or2_1 _8179_ (.A(net327),
    .B(net193),
    .X(_4089_));
 sky130_fd_sc_hd__o211a_1 _8180_ (.A1(net126),
    .A2(net191),
    .B1(_4089_),
    .C1(net214),
    .X(_0548_));
 sky130_fd_sc_hd__or2_1 _8181_ (.A(net359),
    .B(net193),
    .X(_4090_));
 sky130_fd_sc_hd__o211a_1 _8182_ (.A1(net124),
    .A2(net191),
    .B1(_4090_),
    .C1(net214),
    .X(_0549_));
 sky130_fd_sc_hd__or2_1 _8183_ (.A(net377),
    .B(net193),
    .X(_4091_));
 sky130_fd_sc_hd__o211a_1 _8184_ (.A1(net122),
    .A2(net191),
    .B1(_4091_),
    .C1(net213),
    .X(_0550_));
 sky130_fd_sc_hd__or2_1 _8185_ (.A(net391),
    .B(net193),
    .X(_4092_));
 sky130_fd_sc_hd__o211a_1 _8186_ (.A1(net119),
    .A2(net191),
    .B1(_4092_),
    .C1(net213),
    .X(_0551_));
 sky130_fd_sc_hd__or2_1 _8187_ (.A(net395),
    .B(net192),
    .X(_4093_));
 sky130_fd_sc_hd__o211a_1 _8188_ (.A1(net116),
    .A2(net190),
    .B1(_4093_),
    .C1(net212),
    .X(_0552_));
 sky130_fd_sc_hd__or2_1 _8189_ (.A(net357),
    .B(net193),
    .X(_4094_));
 sky130_fd_sc_hd__o211a_1 _8190_ (.A1(net113),
    .A2(net191),
    .B1(_4094_),
    .C1(net213),
    .X(_0553_));
 sky130_fd_sc_hd__or2_1 _8191_ (.A(net397),
    .B(net192),
    .X(_4095_));
 sky130_fd_sc_hd__o211a_1 _8192_ (.A1(net110),
    .A2(net190),
    .B1(_4095_),
    .C1(net211),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _8193_ (.A(net355),
    .B(net192),
    .X(_4096_));
 sky130_fd_sc_hd__o211a_1 _8194_ (.A1(net108),
    .A2(net190),
    .B1(_4096_),
    .C1(net212),
    .X(_0555_));
 sky130_fd_sc_hd__or2_1 _8195_ (.A(net383),
    .B(net192),
    .X(_4097_));
 sky130_fd_sc_hd__o211a_1 _8196_ (.A1(net106),
    .A2(net190),
    .B1(_4097_),
    .C1(net213),
    .X(_0556_));
 sky130_fd_sc_hd__dfxtp_1 _8197_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net403),
    .Q(\ann.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8198_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(\ann.next_state[1] ),
    .Q(\ann.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8199_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0068_),
    .Q(\ann.multiply_FF[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8200_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0069_),
    .Q(\ann.multiply_FF[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8201_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0070_),
    .Q(\ann.multiply_FF[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8202_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0071_),
    .Q(\ann.multiply_FF[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8203_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0072_),
    .Q(\ann.multiply_FF[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8204_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0073_),
    .Q(\ann.multiply_FF[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8205_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0074_),
    .Q(\ann.multiply_FF[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8206_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0075_),
    .Q(\ann.multiply_FF[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8207_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0076_),
    .Q(\ann.multiply_FF[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8208_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0077_),
    .Q(\ann.multiply_FF[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8209_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0078_),
    .Q(\ann.multiply_FF[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8210_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0079_),
    .Q(\ann.multiply_FF[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8211_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0080_),
    .Q(\ann.multiply_FF[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8212_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0081_),
    .Q(\ann.multiply_FF[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8213_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0082_),
    .Q(\ann.multiply_FF[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8214_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0083_),
    .Q(\ann.multiply_FF[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8215_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0084_),
    .Q(\ann.multiply_FF[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8216_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0085_),
    .Q(\ann.multiply_FF[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8217_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0086_),
    .Q(\ann.multiply_FF[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8218_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0087_),
    .Q(\ann.multiply_FF[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8219_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0088_),
    .Q(\ann.multiply_FF[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8220_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0089_),
    .Q(\ann.multiply_FF[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8221_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0090_),
    .Q(\ann.multiply_FF[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8222_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0091_),
    .Q(\ann.multiply_FF[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8223_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0092_),
    .Q(\ann.multiply_FF[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8224_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0093_),
    .Q(\ann.multiply_FF[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8225_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0094_),
    .Q(\ann.multiply_FF[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8226_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0095_),
    .Q(\ann.multiply_FF[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8227_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0096_),
    .Q(\ann.multiply_FF[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8228_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0097_),
    .Q(\ann.multiply_FF[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8229_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0098_),
    .Q(\ann.multiply_FF[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8230_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0099_),
    .Q(\ann.multiply_FF[31] ));
 sky130_fd_sc_hd__dfxtp_4 _8231_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0100_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _8232_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0101_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _8233_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0102_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _8234_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0103_),
    .Q(net35));
 sky130_fd_sc_hd__dlxtn_1 _8235_ (.D(_0032_),
    .GATE_N(net61),
    .Q(\ann.sum[0] ));
 sky130_fd_sc_hd__dlxtn_1 _8236_ (.D(_0043_),
    .GATE_N(net61),
    .Q(\ann.sum[1] ));
 sky130_fd_sc_hd__dlxtn_1 _8237_ (.D(_0054_),
    .GATE_N(net60),
    .Q(\ann.sum[2] ));
 sky130_fd_sc_hd__dlxtn_1 _8238_ (.D(_0057_),
    .GATE_N(net61),
    .Q(\ann.sum[3] ));
 sky130_fd_sc_hd__dlxtn_1 _8239_ (.D(_0058_),
    .GATE_N(net60),
    .Q(\ann.sum[4] ));
 sky130_fd_sc_hd__dlxtn_1 _8240_ (.D(_0059_),
    .GATE_N(net60),
    .Q(\ann.sum[5] ));
 sky130_fd_sc_hd__dlxtn_1 _8241_ (.D(_0060_),
    .GATE_N(_0066_),
    .Q(\ann.sum[6] ));
 sky130_fd_sc_hd__dlxtn_1 _8242_ (.D(_0061_),
    .GATE_N(net61),
    .Q(\ann.sum[7] ));
 sky130_fd_sc_hd__dlxtn_1 _8243_ (.D(_0062_),
    .GATE_N(net61),
    .Q(\ann.sum[8] ));
 sky130_fd_sc_hd__dlxtn_1 _8244_ (.D(_0063_),
    .GATE_N(net61),
    .Q(\ann.sum[9] ));
 sky130_fd_sc_hd__dlxtn_2 _8245_ (.D(_0033_),
    .GATE_N(net61),
    .Q(\ann.sum[10] ));
 sky130_fd_sc_hd__dlxtn_1 _8246_ (.D(_0034_),
    .GATE_N(net61),
    .Q(\ann.sum[11] ));
 sky130_fd_sc_hd__dlxtn_1 _8247_ (.D(_0035_),
    .GATE_N(net61),
    .Q(\ann.sum[12] ));
 sky130_fd_sc_hd__dlxtn_1 _8248_ (.D(_0036_),
    .GATE_N(net61),
    .Q(\ann.sum[13] ));
 sky130_fd_sc_hd__dlxtn_1 _8249_ (.D(_0037_),
    .GATE_N(net61),
    .Q(\ann.sum[14] ));
 sky130_fd_sc_hd__dlxtn_1 _8250_ (.D(_0038_),
    .GATE_N(net61),
    .Q(\ann.sum[15] ));
 sky130_fd_sc_hd__dlxtn_1 _8251_ (.D(_0039_),
    .GATE_N(net61),
    .Q(\ann.sum[16] ));
 sky130_fd_sc_hd__dlxtn_1 _8252_ (.D(_0040_),
    .GATE_N(net60),
    .Q(\ann.sum[17] ));
 sky130_fd_sc_hd__dlxtn_1 _8253_ (.D(_0041_),
    .GATE_N(net60),
    .Q(\ann.sum[18] ));
 sky130_fd_sc_hd__dlxtn_1 _8254_ (.D(_0042_),
    .GATE_N(net60),
    .Q(\ann.sum[19] ));
 sky130_fd_sc_hd__dlxtn_1 _8255_ (.D(_0044_),
    .GATE_N(net60),
    .Q(\ann.sum[20] ));
 sky130_fd_sc_hd__dlxtn_1 _8256_ (.D(_0045_),
    .GATE_N(net60),
    .Q(\ann.sum[21] ));
 sky130_fd_sc_hd__dlxtn_1 _8257_ (.D(_0046_),
    .GATE_N(net60),
    .Q(\ann.sum[22] ));
 sky130_fd_sc_hd__dlxtn_1 _8258_ (.D(_0047_),
    .GATE_N(net60),
    .Q(\ann.sum[23] ));
 sky130_fd_sc_hd__dlxtn_1 _8259_ (.D(_0048_),
    .GATE_N(net60),
    .Q(\ann.sum[24] ));
 sky130_fd_sc_hd__dlxtn_1 _8260_ (.D(_0049_),
    .GATE_N(net60),
    .Q(\ann.sum[25] ));
 sky130_fd_sc_hd__dlxtn_1 _8261_ (.D(_0050_),
    .GATE_N(net60),
    .Q(\ann.sum[26] ));
 sky130_fd_sc_hd__dlxtn_1 _8262_ (.D(_0051_),
    .GATE_N(net60),
    .Q(\ann.sum[27] ));
 sky130_fd_sc_hd__dlxtn_1 _8263_ (.D(_0052_),
    .GATE_N(net60),
    .Q(\ann.sum[28] ));
 sky130_fd_sc_hd__dlxtn_1 _8264_ (.D(_0053_),
    .GATE_N(net60),
    .Q(\ann.sum[29] ));
 sky130_fd_sc_hd__dlxtn_1 _8265_ (.D(_0055_),
    .GATE_N(net61),
    .Q(\ann.sum[30] ));
 sky130_fd_sc_hd__dlxtn_1 _8266_ (.D(_0056_),
    .GATE_N(net61),
    .Q(\ann.sum[31] ));
 sky130_fd_sc_hd__dlxtn_1 _8267_ (.D(_0000_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[0] ));
 sky130_fd_sc_hd__dlxtn_1 _8268_ (.D(_0011_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[1] ));
 sky130_fd_sc_hd__dlxtn_1 _8269_ (.D(_0022_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[2] ));
 sky130_fd_sc_hd__dlxtn_1 _8270_ (.D(_0025_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[3] ));
 sky130_fd_sc_hd__dlxtn_1 _8271_ (.D(_0026_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[4] ));
 sky130_fd_sc_hd__dlxtn_1 _8272_ (.D(_0027_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[5] ));
 sky130_fd_sc_hd__dlxtn_1 _8273_ (.D(_0028_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[6] ));
 sky130_fd_sc_hd__dlxtn_1 _8274_ (.D(_0029_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[7] ));
 sky130_fd_sc_hd__dlxtn_1 _8275_ (.D(_0030_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[8] ));
 sky130_fd_sc_hd__dlxtn_1 _8276_ (.D(_0031_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[9] ));
 sky130_fd_sc_hd__dlxtn_1 _8277_ (.D(_0001_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[10] ));
 sky130_fd_sc_hd__dlxtn_1 _8278_ (.D(_0002_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[11] ));
 sky130_fd_sc_hd__dlxtn_1 _8279_ (.D(_0003_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[12] ));
 sky130_fd_sc_hd__dlxtn_1 _8280_ (.D(_0004_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[13] ));
 sky130_fd_sc_hd__dlxtn_1 _8281_ (.D(_0005_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[14] ));
 sky130_fd_sc_hd__dlxtn_1 _8282_ (.D(_0006_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[15] ));
 sky130_fd_sc_hd__dlxtn_1 _8283_ (.D(_0007_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[16] ));
 sky130_fd_sc_hd__dlxtn_1 _8284_ (.D(_0008_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[17] ));
 sky130_fd_sc_hd__dlxtn_1 _8285_ (.D(_0009_),
    .GATE_N(net92),
    .Q(\ann.multiply_out[18] ));
 sky130_fd_sc_hd__dlxtn_1 _8286_ (.D(_0010_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[19] ));
 sky130_fd_sc_hd__dlxtn_1 _8287_ (.D(_0012_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[20] ));
 sky130_fd_sc_hd__dlxtn_1 _8288_ (.D(_0013_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[21] ));
 sky130_fd_sc_hd__dlxtn_1 _8289_ (.D(_0014_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[22] ));
 sky130_fd_sc_hd__dlxtn_1 _8290_ (.D(_0015_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[23] ));
 sky130_fd_sc_hd__dlxtn_1 _8291_ (.D(_0016_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[24] ));
 sky130_fd_sc_hd__dlxtn_1 _8292_ (.D(_0017_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[25] ));
 sky130_fd_sc_hd__dlxtn_1 _8293_ (.D(_0018_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[26] ));
 sky130_fd_sc_hd__dlxtn_1 _8294_ (.D(_0019_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[27] ));
 sky130_fd_sc_hd__dlxtn_1 _8295_ (.D(_0020_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[28] ));
 sky130_fd_sc_hd__dlxtn_1 _8296_ (.D(_0021_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[29] ));
 sky130_fd_sc_hd__dlxtn_1 _8297_ (.D(_0023_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[30] ));
 sky130_fd_sc_hd__dlxtn_1 _8298_ (.D(_0024_),
    .GATE_N(net91),
    .Q(\ann.multiply_out[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8299_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net354),
    .Q(\ann.temp[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8300_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net366),
    .Q(\ann.temp[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8301_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net344),
    .Q(\ann.temp[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8302_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net350),
    .Q(\ann.temp[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8303_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net352),
    .Q(\ann.temp[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8304_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net330),
    .Q(\ann.temp[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8305_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net380),
    .Q(\ann.temp[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8306_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net334),
    .Q(\ann.temp[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8307_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0112_),
    .Q(\ann.temp[8] ));
 sky130_fd_sc_hd__dfxtp_2 _8308_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0113_),
    .Q(\ann.temp[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8309_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0114_),
    .Q(\ann.temp[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8310_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0115_),
    .Q(\ann.temp[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8311_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net340),
    .Q(\ann.temp[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8312_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net316),
    .Q(\ann.temp[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8313_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net314),
    .Q(\ann.temp[14] ));
 sky130_fd_sc_hd__dfxtp_4 _8314_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0119_),
    .Q(\ann.temp[15] ));
 sky130_fd_sc_hd__dfxtp_2 _8315_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0120_),
    .Q(\ann.temp[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8316_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0121_),
    .Q(\ann.temp[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8317_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0122_),
    .Q(\ann.temp[18] ));
 sky130_fd_sc_hd__dfxtp_4 _8318_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0123_),
    .Q(\ann.temp[19] ));
 sky130_fd_sc_hd__dfxtp_2 _8319_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0124_),
    .Q(\ann.temp[20] ));
 sky130_fd_sc_hd__dfxtp_2 _8320_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0125_),
    .Q(\ann.temp[21] ));
 sky130_fd_sc_hd__dfxtp_2 _8321_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0126_),
    .Q(\ann.temp[22] ));
 sky130_fd_sc_hd__dfxtp_2 _8322_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0127_),
    .Q(\ann.temp[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8323_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0128_),
    .Q(\ann.temp[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8324_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0129_),
    .Q(\ann.temp[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8325_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0130_),
    .Q(\ann.temp[26] ));
 sky130_fd_sc_hd__dfxtp_4 _8326_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0131_),
    .Q(\ann.temp[27] ));
 sky130_fd_sc_hd__dfxtp_4 _8327_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0132_),
    .Q(\ann.temp[28] ));
 sky130_fd_sc_hd__dfxtp_4 _8328_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0133_),
    .Q(\ann.temp[29] ));
 sky130_fd_sc_hd__dfxtp_2 _8329_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0134_),
    .Q(\ann.temp[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8330_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net288),
    .Q(\ann.ReLU_out[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8331_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net264),
    .Q(\ann.ReLU_out[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8332_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net284),
    .Q(\ann.ReLU_out[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8333_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net304),
    .Q(\ann.ReLU_out[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8334_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net296),
    .Q(\ann.ReLU_out[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8335_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net298),
    .Q(\ann.ReLU_out[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8336_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net292),
    .Q(\ann.ReLU_out[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8337_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net278),
    .Q(\ann.ReLU_out[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8338_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net306),
    .Q(\ann.ReLU_out[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8339_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net262),
    .Q(\ann.ReLU_out[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8340_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net276),
    .Q(\ann.ReLU_out[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8341_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net302),
    .Q(\ann.ReLU_out[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8342_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net270),
    .Q(\ann.ReLU_out[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8343_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net266),
    .Q(\ann.ReLU_out[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8344_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net260),
    .Q(\ann.ReLU_out[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8345_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net318),
    .Q(\ann.ReLU_out[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8346_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net280),
    .Q(\ann.ReLU_out[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8347_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net272),
    .Q(\ann.ReLU_out[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8348_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net268),
    .Q(\ann.ReLU_out[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8349_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net308),
    .Q(\ann.ReLU_out[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8350_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net286),
    .Q(\ann.ReLU_out[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8351_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net256),
    .Q(\ann.ReLU_out[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8352_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net300),
    .Q(\ann.ReLU_out[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8353_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net282),
    .Q(\ann.ReLU_out[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8354_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net290),
    .Q(\ann.ReLU_out[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8355_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net310),
    .Q(\ann.ReLU_out[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8356_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net320),
    .Q(\ann.ReLU_out[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8357_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net294),
    .Q(\ann.ReLU_out[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8358_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net312),
    .Q(\ann.ReLU_out[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8359_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net274),
    .Q(\ann.ReLU_out[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8360_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net258),
    .Q(\ann.ReLU_out[0][30] ));
 sky130_fd_sc_hd__dlxtn_1 _8361_ (.D(_0558_),
    .GATE_N(_0065_),
    .Q(\ann.add_enable ));
 sky130_fd_sc_hd__dfxtp_1 _8362_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net324),
    .Q(\ann.ReLU_out[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8363_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0167_),
    .Q(\ann.ReLU_out[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8364_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0168_),
    .Q(\ann.ReLU_out[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8365_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0169_),
    .Q(\ann.ReLU_out[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8366_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0170_),
    .Q(\ann.ReLU_out[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8367_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0171_),
    .Q(\ann.ReLU_out[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8368_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0172_),
    .Q(\ann.ReLU_out[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8369_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0173_),
    .Q(\ann.ReLU_out[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8370_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0174_),
    .Q(\ann.ReLU_out[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8371_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0175_),
    .Q(\ann.ReLU_out[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8372_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0176_),
    .Q(\ann.ReLU_out[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8373_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0177_),
    .Q(\ann.ReLU_out[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8374_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0178_),
    .Q(\ann.ReLU_out[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8375_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0179_),
    .Q(\ann.ReLU_out[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8376_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0180_),
    .Q(\ann.ReLU_out[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8377_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0181_),
    .Q(\ann.ReLU_out[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8378_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0182_),
    .Q(\ann.ReLU_out[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8379_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0183_),
    .Q(\ann.ReLU_out[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8380_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0184_),
    .Q(\ann.ReLU_out[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8381_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0185_),
    .Q(\ann.ReLU_out[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8382_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0186_),
    .Q(\ann.ReLU_out[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8383_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0187_),
    .Q(\ann.ReLU_out[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _8384_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0188_),
    .Q(\ann.ReLU_out[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8385_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0189_),
    .Q(\ann.ReLU_out[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8386_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0190_),
    .Q(\ann.ReLU_out[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8387_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0191_),
    .Q(\ann.ReLU_out[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8388_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0192_),
    .Q(\ann.ReLU_out[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8389_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0193_),
    .Q(\ann.ReLU_out[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8390_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0194_),
    .Q(\ann.ReLU_out[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8391_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0195_),
    .Q(\ann.ReLU_out[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8392_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0196_),
    .Q(\ann.ReLU_out[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8393_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net326),
    .Q(\ann.ReLU_out[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8394_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0198_),
    .Q(\ann.ReLU_out[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8395_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0199_),
    .Q(\ann.ReLU_out[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8396_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0200_),
    .Q(\ann.ReLU_out[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8397_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0201_),
    .Q(\ann.ReLU_out[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8398_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0202_),
    .Q(\ann.ReLU_out[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8399_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0203_),
    .Q(\ann.ReLU_out[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8400_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0204_),
    .Q(\ann.ReLU_out[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8401_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0205_),
    .Q(\ann.ReLU_out[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8402_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0206_),
    .Q(\ann.ReLU_out[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8403_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0207_),
    .Q(\ann.ReLU_out[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8404_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0208_),
    .Q(\ann.ReLU_out[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8405_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0209_),
    .Q(\ann.ReLU_out[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8406_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0210_),
    .Q(\ann.ReLU_out[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8407_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0211_),
    .Q(\ann.ReLU_out[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8408_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0212_),
    .Q(\ann.ReLU_out[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8409_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net401),
    .Q(\ann.ReLU_out[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8410_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net416),
    .Q(\ann.ReLU_out[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8411_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0215_),
    .Q(\ann.ReLU_out[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8412_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0216_),
    .Q(\ann.ReLU_out[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8413_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0217_),
    .Q(\ann.ReLU_out[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8414_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0218_),
    .Q(\ann.ReLU_out[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8415_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0219_),
    .Q(\ann.ReLU_out[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8416_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0220_),
    .Q(\ann.ReLU_out[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8417_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0221_),
    .Q(\ann.ReLU_out[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8418_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0222_),
    .Q(\ann.ReLU_out[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8419_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0223_),
    .Q(\ann.ReLU_out[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8420_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0224_),
    .Q(\ann.ReLU_out[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8421_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0225_),
    .Q(\ann.ReLU_out[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8422_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0226_),
    .Q(\ann.ReLU_out[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8423_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0227_),
    .Q(\ann.ReLU_out[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8424_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net342),
    .Q(\ann.ReLU_out[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8425_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0229_),
    .Q(\ann.ReLU_out[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8426_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0230_),
    .Q(\ann.ReLU_out[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8427_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0231_),
    .Q(\ann.ReLU_out[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8428_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0232_),
    .Q(\ann.ReLU_out[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8429_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0233_),
    .Q(\ann.ReLU_out[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8430_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0234_),
    .Q(\ann.ReLU_out[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8431_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0235_),
    .Q(\ann.ReLU_out[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8432_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0236_),
    .Q(\ann.ReLU_out[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8433_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0237_),
    .Q(\ann.ReLU_out[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8434_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0238_),
    .Q(\ann.ReLU_out[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8435_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0239_),
    .Q(\ann.ReLU_out[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8436_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0240_),
    .Q(\ann.ReLU_out[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8437_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0241_),
    .Q(\ann.ReLU_out[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8438_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0242_),
    .Q(\ann.ReLU_out[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8439_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0243_),
    .Q(\ann.ReLU_out[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8440_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0244_),
    .Q(\ann.ReLU_out[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8441_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0245_),
    .Q(\ann.ReLU_out[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8442_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0246_),
    .Q(\ann.ReLU_out[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8443_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0247_),
    .Q(\ann.ReLU_out[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8444_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0248_),
    .Q(\ann.ReLU_out[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8445_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0249_),
    .Q(\ann.ReLU_out[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8446_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0250_),
    .Q(\ann.ReLU_out[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8447_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0251_),
    .Q(\ann.ReLU_out[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8448_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0252_),
    .Q(\ann.ReLU_out[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8449_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0253_),
    .Q(\ann.ReLU_out[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8450_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0254_),
    .Q(\ann.ReLU_out[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8451_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0255_),
    .Q(\ann.ReLU_out[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8452_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0256_),
    .Q(\ann.ReLU_out[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8453_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0257_),
    .Q(\ann.ReLU_out[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8454_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net390),
    .Q(\ann.ReLU_out[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8455_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net388),
    .Q(\ann.ReLU_out[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8456_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0260_),
    .Q(\ann.ReLU_out[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8457_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0261_),
    .Q(\ann.ReLU_out[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8458_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0262_),
    .Q(\ann.ReLU_out[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8459_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0263_),
    .Q(\ann.ReLU_out[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8460_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0264_),
    .Q(\ann.ReLU_out[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8461_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0265_),
    .Q(\ann.ReLU_out[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8462_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0266_),
    .Q(\ann.ReLU_out[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8463_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0267_),
    .Q(\ann.ReLU_out[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8464_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0268_),
    .Q(\ann.ReLU_out[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8465_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0269_),
    .Q(\ann.ReLU_out[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8466_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0270_),
    .Q(\ann.ReLU_out[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8467_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0271_),
    .Q(\ann.ReLU_out[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8468_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0272_),
    .Q(\ann.ReLU_out[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8469_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0273_),
    .Q(\ann.ReLU_out[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8470_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0274_),
    .Q(\ann.ReLU_out[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8471_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0275_),
    .Q(\ann.ReLU_out[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8472_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0276_),
    .Q(\ann.ReLU_out[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8473_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0277_),
    .Q(\ann.ReLU_out[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8474_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0278_),
    .Q(\ann.ReLU_out[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8475_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0279_),
    .Q(\ann.ReLU_out[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8476_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0280_),
    .Q(\ann.ReLU_out[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8477_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0281_),
    .Q(\ann.ReLU_out[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8478_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0282_),
    .Q(\ann.ReLU_out[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8479_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0283_),
    .Q(\ann.ReLU_out[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8480_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0284_),
    .Q(\ann.ReLU_out[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8481_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0285_),
    .Q(\ann.ReLU_out[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8482_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0286_),
    .Q(\ann.ReLU_out[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8483_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0287_),
    .Q(\ann.ReLU_out[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8484_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0288_),
    .Q(\ann.ReLU_out[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8485_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0289_),
    .Q(\ann.ReLU_out[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8486_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net348),
    .Q(\ann.ReLU_out[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8487_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0291_),
    .Q(\ann.ReLU_out[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8488_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0292_),
    .Q(\ann.ReLU_out[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8489_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0293_),
    .Q(\ann.ReLU_out[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8490_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0294_),
    .Q(\ann.ReLU_out[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8491_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0295_),
    .Q(\ann.ReLU_out[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8492_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net467),
    .Q(\ann.ReLU_out[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8493_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0297_),
    .Q(\ann.ReLU_out[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8494_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0298_),
    .Q(\ann.ReLU_out[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8495_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0299_),
    .Q(\ann.ReLU_out[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8496_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0300_),
    .Q(\ann.ReLU_out[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8497_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0301_),
    .Q(\ann.ReLU_out[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8498_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0302_),
    .Q(\ann.ReLU_out[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8499_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0303_),
    .Q(\ann.ReLU_out[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8500_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0304_),
    .Q(\ann.ReLU_out[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8501_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0305_),
    .Q(\ann.ReLU_out[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8502_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0306_),
    .Q(\ann.ReLU_out[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8503_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0307_),
    .Q(\ann.ReLU_out[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8504_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0308_),
    .Q(\ann.ReLU_out[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8505_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0309_),
    .Q(\ann.ReLU_out[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8506_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0310_),
    .Q(\ann.ReLU_out[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8507_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0311_),
    .Q(\ann.ReLU_out[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8508_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0312_),
    .Q(\ann.ReLU_out[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8509_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0313_),
    .Q(\ann.ReLU_out[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8510_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0314_),
    .Q(\ann.ReLU_out[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8511_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0315_),
    .Q(\ann.ReLU_out[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8512_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0316_),
    .Q(\ann.ReLU_out[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8513_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0317_),
    .Q(\ann.ReLU_out[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8514_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0318_),
    .Q(\ann.ReLU_out[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8515_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net405),
    .Q(\ann.ReLU_out[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8516_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0320_),
    .Q(\ann.ReLU_out[5][30] ));
 sky130_fd_sc_hd__dlxtn_1 _8517_ (.D(_0557_),
    .GATE_N(net223),
    .Q(\ann.ldX ));
 sky130_fd_sc_hd__conb_1 _8517__223 (.LO(net223));
 sky130_fd_sc_hd__dfxtp_1 _8518_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net386),
    .Q(\ann.ReLU_out[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8519_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0322_),
    .Q(\ann.ReLU_out[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8520_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0323_),
    .Q(\ann.ReLU_out[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8521_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0324_),
    .Q(\ann.ReLU_out[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8522_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0325_),
    .Q(\ann.ReLU_out[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8523_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0326_),
    .Q(\ann.ReLU_out[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8524_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0327_),
    .Q(\ann.ReLU_out[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8525_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0328_),
    .Q(\ann.ReLU_out[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8526_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net338),
    .Q(\ann.ReLU_out[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8527_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0330_),
    .Q(\ann.ReLU_out[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8528_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0331_),
    .Q(\ann.ReLU_out[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8529_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0332_),
    .Q(\ann.ReLU_out[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8530_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net409),
    .Q(\ann.ReLU_out[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8531_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0334_),
    .Q(\ann.ReLU_out[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8532_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0335_),
    .Q(\ann.ReLU_out[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8533_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0336_),
    .Q(\ann.ReLU_out[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8534_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net370),
    .Q(\ann.ReLU_out[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8535_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net336),
    .Q(\ann.ReLU_out[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8536_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0339_),
    .Q(\ann.ReLU_out[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8537_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0340_),
    .Q(\ann.ReLU_out[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8538_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0341_),
    .Q(\ann.ReLU_out[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8539_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0342_),
    .Q(\ann.ReLU_out[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8540_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0343_),
    .Q(\ann.ReLU_out[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8541_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0344_),
    .Q(\ann.ReLU_out[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8542_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0345_),
    .Q(\ann.ReLU_out[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8543_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0346_),
    .Q(\ann.ReLU_out[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8544_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0347_),
    .Q(\ann.ReLU_out[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8545_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0348_),
    .Q(\ann.ReLU_out[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8546_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0349_),
    .Q(\ann.ReLU_out[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8547_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0350_),
    .Q(\ann.ReLU_out[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8548_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net322),
    .Q(\ann.ReLU_out[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8549_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net368),
    .Q(\ann.ReLU_out[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8550_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0353_),
    .Q(\ann.ReLU_out[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8551_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0354_),
    .Q(\ann.ReLU_out[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8552_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0355_),
    .Q(\ann.ReLU_out[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8553_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0356_),
    .Q(\ann.ReLU_out[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8554_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0357_),
    .Q(\ann.ReLU_out[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8555_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0358_),
    .Q(\ann.ReLU_out[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8556_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0359_),
    .Q(\ann.ReLU_out[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8557_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0360_),
    .Q(\ann.ReLU_out[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8558_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0361_),
    .Q(\ann.ReLU_out[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8559_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0362_),
    .Q(\ann.ReLU_out[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8560_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0363_),
    .Q(\ann.ReLU_out[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8561_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0364_),
    .Q(\ann.ReLU_out[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8562_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0365_),
    .Q(\ann.ReLU_out[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8563_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0366_),
    .Q(\ann.ReLU_out[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8564_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0367_),
    .Q(\ann.ReLU_out[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8565_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0368_),
    .Q(\ann.ReLU_out[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8566_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0369_),
    .Q(\ann.ReLU_out[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8567_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0370_),
    .Q(\ann.ReLU_out[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8568_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0371_),
    .Q(\ann.ReLU_out[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8569_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0372_),
    .Q(\ann.ReLU_out[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8570_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0373_),
    .Q(\ann.ReLU_out[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8571_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0374_),
    .Q(\ann.ReLU_out[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8572_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0375_),
    .Q(\ann.ReLU_out[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8573_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0376_),
    .Q(\ann.ReLU_out[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8574_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0377_),
    .Q(\ann.ReLU_out[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8575_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0378_),
    .Q(\ann.ReLU_out[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8576_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0379_),
    .Q(\ann.ReLU_out[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8577_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0380_),
    .Q(\ann.ReLU_out[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8578_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0381_),
    .Q(\ann.ReLU_out[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8579_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0382_),
    .Q(\ann.ReLU_out[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8580_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net382),
    .Q(\ann.ReLU_out[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8581_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0384_),
    .Q(\ann.ReLU_out[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8582_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0385_),
    .Q(\ann.ReLU_out[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8583_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0386_),
    .Q(\ann.ReLU_out[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8584_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0387_),
    .Q(\ann.ReLU_out[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8585_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0388_),
    .Q(\ann.ReLU_out[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8586_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0389_),
    .Q(\ann.ReLU_out[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8587_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0390_),
    .Q(\ann.ReLU_out[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8588_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0391_),
    .Q(\ann.ReLU_out[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8589_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0392_),
    .Q(\ann.ReLU_out[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8590_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0393_),
    .Q(\ann.ReLU_out[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8591_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0394_),
    .Q(\ann.ReLU_out[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8592_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0395_),
    .Q(\ann.ReLU_out[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8593_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0396_),
    .Q(\ann.ReLU_out[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8594_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0397_),
    .Q(\ann.ReLU_out[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8595_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0398_),
    .Q(\ann.ReLU_out[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8596_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0399_),
    .Q(\ann.ReLU_out[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8597_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0400_),
    .Q(\ann.ReLU_out[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8598_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0401_),
    .Q(\ann.ReLU_out[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8599_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0402_),
    .Q(\ann.ReLU_out[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8600_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0403_),
    .Q(\ann.ReLU_out[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8601_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0404_),
    .Q(\ann.ReLU_out[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8602_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0405_),
    .Q(\ann.ReLU_out[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8603_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0406_),
    .Q(\ann.ReLU_out[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8604_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0407_),
    .Q(\ann.ReLU_out[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8605_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0408_),
    .Q(\ann.ReLU_out[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8606_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0409_),
    .Q(\ann.ReLU_out[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8607_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0410_),
    .Q(\ann.ReLU_out[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8608_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0411_),
    .Q(\ann.ReLU_out[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8609_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0412_),
    .Q(\ann.ReLU_out[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8610_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0413_),
    .Q(\ann.ReLU_out[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8611_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0414_),
    .Q(\ann.X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8612_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0415_),
    .Q(\ann.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8613_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0416_),
    .Q(\ann.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8614_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0417_),
    .Q(\ann.X[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8615_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0418_),
    .Q(\ann.X[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8616_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0419_),
    .Q(\ann.X[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8617_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0420_),
    .Q(\ann.X[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8618_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0421_),
    .Q(\ann.X[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8619_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0422_),
    .Q(\ann.X[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8620_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0423_),
    .Q(\ann.X[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8621_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0424_),
    .Q(\ann.X[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8622_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0425_),
    .Q(\ann.X[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8623_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0426_),
    .Q(\ann.X[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8624_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0427_),
    .Q(\ann.X[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8625_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0428_),
    .Q(\ann.X[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8626_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0429_),
    .Q(\ann.X[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8627_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0430_),
    .Q(\ann.X[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8628_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0431_),
    .Q(\ann.X[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8629_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0432_),
    .Q(\ann.X[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8630_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0433_),
    .Q(\ann.X[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8631_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0434_),
    .Q(\ann.X[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8632_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0435_),
    .Q(\ann.X[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8633_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0436_),
    .Q(\ann.X[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8634_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0437_),
    .Q(\ann.X[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8635_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0438_),
    .Q(\ann.X[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8636_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0439_),
    .Q(\ann.X[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8637_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0440_),
    .Q(\ann.X[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8638_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0441_),
    .Q(\ann.X[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8639_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0442_),
    .Q(\ann.X[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8640_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0443_),
    .Q(\ann.X[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8641_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0444_),
    .Q(\ann.X[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8642_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0445_),
    .Q(\ann.X[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8643_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net394),
    .Q(\ann.ReLU_out[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8644_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0447_),
    .Q(\ann.ReLU_out[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8645_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0448_),
    .Q(\ann.ReLU_out[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8646_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0449_),
    .Q(\ann.ReLU_out[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8647_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0450_),
    .Q(\ann.ReLU_out[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8648_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0451_),
    .Q(\ann.ReLU_out[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8649_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0452_),
    .Q(\ann.ReLU_out[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8650_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0453_),
    .Q(\ann.ReLU_out[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8651_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0454_),
    .Q(\ann.ReLU_out[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8652_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0455_),
    .Q(\ann.ReLU_out[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8653_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0456_),
    .Q(\ann.ReLU_out[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8654_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0457_),
    .Q(\ann.ReLU_out[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8655_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0458_),
    .Q(\ann.ReLU_out[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8656_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0459_),
    .Q(\ann.ReLU_out[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8657_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0460_),
    .Q(\ann.ReLU_out[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8658_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0461_),
    .Q(\ann.ReLU_out[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8659_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0462_),
    .Q(\ann.ReLU_out[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _8660_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0463_),
    .Q(\ann.ReLU_out[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _8661_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0464_),
    .Q(\ann.ReLU_out[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _8662_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0465_),
    .Q(\ann.ReLU_out[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _8663_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0466_),
    .Q(\ann.ReLU_out[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _8664_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0467_),
    .Q(\ann.ReLU_out[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _8665_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0468_),
    .Q(\ann.ReLU_out[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _8666_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0469_),
    .Q(\ann.ReLU_out[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _8667_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0470_),
    .Q(\ann.ReLU_out[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _8668_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0471_),
    .Q(\ann.ReLU_out[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _8669_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0472_),
    .Q(\ann.ReLU_out[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _8670_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0473_),
    .Q(\ann.ReLU_out[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _8671_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0474_),
    .Q(\ann.ReLU_out[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _8672_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0475_),
    .Q(\ann.ReLU_out[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _8673_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0476_),
    .Q(\ann.ReLU_out[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _8674_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0477_),
    .Q(\ann.bias[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8675_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0478_),
    .Q(\ann.bias[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8676_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0479_),
    .Q(\ann.bias[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8677_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0480_),
    .Q(\ann.bias[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8678_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0481_),
    .Q(\ann.bias[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8679_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0482_),
    .Q(\ann.bias[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8680_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0483_),
    .Q(\ann.bias[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8681_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0484_),
    .Q(\ann.bias[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8682_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0485_),
    .Q(\ann.bias[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8683_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0486_),
    .Q(\ann.bias[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8684_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0487_),
    .Q(\ann.bias[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8685_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0488_),
    .Q(\ann.bias[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8686_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0489_),
    .Q(\ann.bias[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8687_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0490_),
    .Q(\ann.bias[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8688_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0491_),
    .Q(\ann.bias[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8689_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0492_),
    .Q(\ann.bias[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8690_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0493_),
    .Q(\ann.bias[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8691_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0494_),
    .Q(\ann.bias[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8692_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0495_),
    .Q(\ann.bias[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8693_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0496_),
    .Q(\ann.bias[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8694_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0497_),
    .Q(\ann.bias[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8695_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0498_),
    .Q(\ann.bias[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8696_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0499_),
    .Q(\ann.bias[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8697_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0500_),
    .Q(\ann.bias[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8698_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0501_),
    .Q(\ann.bias[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8699_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0502_),
    .Q(\ann.bias[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8700_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0503_),
    .Q(\ann.bias[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8701_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0504_),
    .Q(\ann.bias[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8702_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0505_),
    .Q(\ann.bias[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8703_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0506_),
    .Q(\ann.bias[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8704_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0507_),
    .Q(\ann.bias[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8705_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0508_),
    .Q(\ann.bias[15] ));
 sky130_fd_sc_hd__dfxtp_2 _8706_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net29),
    .Q(\ann.weight[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8707_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net30),
    .Q(\ann.weight[1] ));
 sky130_fd_sc_hd__dfxtp_4 _8708_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1),
    .Q(\ann.weight[2] ));
 sky130_fd_sc_hd__dfxtp_4 _8709_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net2),
    .Q(\ann.weight[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8710_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net3),
    .Q(\ann.weight[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8711_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net4),
    .Q(\ann.weight[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8712_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net5),
    .Q(\ann.weight[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8713_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net6),
    .Q(\ann.weight[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8714_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net7),
    .Q(\ann.weight[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8715_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net8),
    .Q(\ann.weight[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8716_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net9),
    .Q(\ann.weight[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8717_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net10),
    .Q(\ann.weight[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8718_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net11),
    .Q(\ann.weight[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8719_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net12),
    .Q(\ann.weight[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8720_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net13),
    .Q(\ann.weight[14] ));
 sky130_fd_sc_hd__dfxtp_2 _8721_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net14),
    .Q(\ann.weight[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8722_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0509_),
    .Q(\ann.in_ff[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8723_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0510_),
    .Q(\ann.in_ff[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8724_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0511_),
    .Q(\ann.in_ff[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8725_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0512_),
    .Q(\ann.in_ff[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8726_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0513_),
    .Q(\ann.in_ff[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8727_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0514_),
    .Q(\ann.in_ff[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8728_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0515_),
    .Q(\ann.in_ff[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8729_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0516_),
    .Q(\ann.in_ff[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8730_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0517_),
    .Q(\ann.in_ff[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8731_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0518_),
    .Q(\ann.in_ff[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8732_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0519_),
    .Q(\ann.in_ff[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8733_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0520_),
    .Q(\ann.in_ff[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8734_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0521_),
    .Q(\ann.in_ff[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8735_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0522_),
    .Q(\ann.in_ff[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8736_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0523_),
    .Q(\ann.in_ff[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8737_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0524_),
    .Q(\ann.in_ff[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8738_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net332),
    .Q(\ann.in_ff[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8739_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net346),
    .Q(\ann.in_ff[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8740_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net372),
    .Q(\ann.in_ff[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8741_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net374),
    .Q(\ann.in_ff[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8742_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net362),
    .Q(\ann.in_ff[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8743_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net364),
    .Q(\ann.in_ff[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8744_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net376),
    .Q(\ann.in_ff[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8745_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net328),
    .Q(\ann.in_ff[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8746_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net360),
    .Q(\ann.in_ff[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8747_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net378),
    .Q(\ann.in_ff[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8748_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net392),
    .Q(\ann.in_ff[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8749_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net396),
    .Q(\ann.in_ff[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8750_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net358),
    .Q(\ann.in_ff[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8751_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net398),
    .Q(\ann.in_ff[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8752_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net356),
    .Q(\ann.in_ff[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8753_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net384),
    .Q(\ann.in_ff[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8754_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0541_),
    .Q(\ann.in_ff[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8755_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0542_),
    .Q(\ann.in_ff[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8756_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0543_),
    .Q(\ann.in_ff[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8757_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0544_),
    .Q(\ann.in_ff[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8758_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0545_),
    .Q(\ann.in_ff[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8759_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0546_),
    .Q(\ann.in_ff[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _8760_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0547_),
    .Q(\ann.in_ff[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _8761_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0548_),
    .Q(\ann.in_ff[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _8762_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0549_),
    .Q(\ann.in_ff[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8763_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0550_),
    .Q(\ann.in_ff[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8764_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0551_),
    .Q(\ann.in_ff[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8765_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0552_),
    .Q(\ann.in_ff[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8766_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0553_),
    .Q(\ann.in_ff[2][12] ));
 sky130_fd_sc_hd__dfxtp_4 _8767_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0554_),
    .Q(\ann.in_ff[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _8768_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0555_),
    .Q(\ann.in_ff[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8769_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0556_),
    .Q(\ann.in_ff[2][15] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(_0649_),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(_0648_),
    .X(net101));
 sky130_fd_sc_hd__buf_4 fanout102 (.A(_0647_),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(_0646_),
    .X(net103));
 sky130_fd_sc_hd__buf_4 fanout104 (.A(_0567_),
    .X(net104));
 sky130_fd_sc_hd__buf_4 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net654),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_8 fanout108 (.A(net662),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(\ann.in_ff[2][13] ),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout110 (.A(net661),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net611),
    .X(net113));
 sky130_fd_sc_hd__buf_4 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net649),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net668),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net660),
    .X(net122));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_8 fanout124 (.A(net642),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(net619),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_8 fanout128 (.A(net630),
    .X(net128));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net131),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net635),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net134),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net625),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net137),
    .X(net135));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net653),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 fanout138 (.A(net140),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net652),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net457),
    .X(net143));
 sky130_fd_sc_hd__buf_6 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net584),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_8 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(\ann.weight[15] ),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(\ann.weight[15] ),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(\ann.weight[14] ),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(\ann.weight[14] ),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(\ann.weight[13] ),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net155),
    .X(net153));
 sky130_fd_sc_hd__buf_2 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_4 fanout155 (.A(\ann.weight[12] ),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(\ann.weight[11] ),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(\ann.weight[10] ),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(\ann.weight[9] ),
    .X(net163));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_8 fanout165 (.A(\ann.weight[8] ),
    .X(net165));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(\ann.weight[7] ),
    .X(net167));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(\ann.weight[6] ),
    .X(net168));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(\ann.weight[6] ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_8 fanout171 (.A(\ann.weight[5] ),
    .X(net171));
 sky130_fd_sc_hd__buf_2 fanout172 (.A(\ann.weight[5] ),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(\ann.weight[4] ),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(\ann.weight[3] ),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(\ann.weight[3] ),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(\ann.weight[2] ),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(\ann.weight[1] ),
    .X(net179));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_6 fanout181 (.A(\ann.weight[0] ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_8 fanout182 (.A(net773),
    .X(net182));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(\ann.temp[25] ),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(\ann.temp[24] ),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_8 fanout185 (.A(\ann.temp[23] ),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(net785),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net782),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net765),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net758),
    .X(net189));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(_4065_),
    .X(net190));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(_4065_),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(_4064_),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(_4064_),
    .X(net193));
 sky130_fd_sc_hd__buf_6 fanout194 (.A(_0709_),
    .X(net194));
 sky130_fd_sc_hd__buf_4 fanout195 (.A(_0709_),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net209),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net209),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(net209),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net204),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(net209),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_2 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_2 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 fanout209 (.A(_0708_),
    .X(net209));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(net215),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net215),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(_0564_),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net27),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(net25),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_8 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_6 fanout37 (.A(_3507_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_8 fanout39 (.A(_3142_),
    .X(net39));
 sky130_fd_sc_hd__buf_6 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_8 fanout41 (.A(_3629_),
    .X(net41));
 sky130_fd_sc_hd__buf_6 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_6 fanout43 (.A(_3566_),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_8 fanout44 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_6 fanout46 (.A(_3324_),
    .X(net46));
 sky130_fd_sc_hd__buf_6 fanout47 (.A(net49),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_6 fanout49 (.A(_3266_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 fanout50 (.A(net52),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_6 fanout52 (.A(_3204_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_6 fanout54 (.A(_3444_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(_3384_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(\ann.sum[31] ),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(_0066_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(_0566_),
    .X(net63));
 sky130_fd_sc_hd__buf_6 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_8 fanout65 (.A(\ann.ldX ),
    .X(net65));
 sky130_fd_sc_hd__buf_4 fanout66 (.A(net68),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(\ann.add_enable ),
    .X(net68));
 sky130_fd_sc_hd__buf_6 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_6 fanout70 (.A(_3999_),
    .X(net70));
 sky130_fd_sc_hd__buf_6 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_8 fanout72 (.A(_3964_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_8 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__buf_6 fanout74 (.A(_3963_),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__buf_8 fanout76 (.A(_3962_),
    .X(net76));
 sky130_fd_sc_hd__buf_6 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_6 fanout78 (.A(_3960_),
    .X(net78));
 sky130_fd_sc_hd__buf_6 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__buf_8 fanout80 (.A(_3966_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_8 fanout81 (.A(_3958_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_8 fanout82 (.A(_3958_),
    .X(net82));
 sky130_fd_sc_hd__buf_6 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_8 fanout84 (.A(_3957_),
    .X(net84));
 sky130_fd_sc_hd__buf_6 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(_3956_),
    .X(net86));
 sky130_fd_sc_hd__buf_6 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_8 fanout88 (.A(_3924_),
    .X(net88));
 sky130_fd_sc_hd__buf_6 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(_3637_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(_0067_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 fanout92 (.A(_0067_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 fanout93 (.A(_0660_),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(_0659_),
    .X(net94));
 sky130_fd_sc_hd__buf_4 fanout95 (.A(_0658_),
    .X(net95));
 sky130_fd_sc_hd__buf_4 fanout96 (.A(_0657_),
    .X(net96));
 sky130_fd_sc_hd__buf_4 fanout97 (.A(_0656_),
    .X(net97));
 sky130_fd_sc_hd__buf_4 fanout98 (.A(_0655_),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(_0654_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\ann.ReLU_out[0][21] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0136_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0104_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\ann.in_ff[1][14] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0539_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\ann.in_ff[1][12] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0537_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\ann.in_ff[1][8] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0533_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\ann.in_ff[1][4] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0529_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\ann.in_ff[1][5] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\ann.ReLU_out[0][13] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0530_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\ann.temp[1] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0105_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\ann.ReLU_out[7][0] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0352_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\ann.ReLU_out[6][16] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0337_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\ann.in_ff[1][2] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0527_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\ann.in_ff[1][3] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0148_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0528_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\ann.in_ff[1][6] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0531_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\ann.in_ff[1][9] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0534_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\ann.temp[6] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0110_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\ann.ReLU_out[8][0] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0383_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\ann.in_ff[1][15] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\ann.ReLU_out[0][18] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0540_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\ann.ReLU_out[6][0] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0321_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\ann.ReLU_out[4][0] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0259_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\ann.ReLU_out[3][30] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0258_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\ann.in_ff[1][10] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0535_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\ann.ReLU_out[9][0] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0153_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0446_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\ann.in_ff[1][11] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0536_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\ann.in_ff[1][13] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0538_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\ann.ReLU_out[6][22] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\ann.ReLU_out[2][16] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0213_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\ann.state[1] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\ann.next_state[0] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\ann.ReLU_out[0][12] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\ann.ReLU_out[5][29] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0319_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\ann.ReLU_out[9][17] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\ann.ReLU_out[3][8] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\ann.ReLU_out[6][12] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0333_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\ann.ReLU_out[1][16] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\ann.ReLU_out[8][24] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\ann.ReLU_out[4][16] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\ann.ReLU_out[3][24] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0147_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\ann.ReLU_out[2][29] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\ann.ReLU_out[2][17] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0214_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\ann.ReLU_out[8][1] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\ann.ReLU_out[8][23] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\ann.ReLU_out[1][18] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\ann.ReLU_out[1][8] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\ann.ReLU_out[6][10] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\ann.ReLU_out[5][22] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\ann.ReLU_out[4][8] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\ann.ReLU_out[0][17] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\ann.ReLU_out[7][23] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\ann.ReLU_out[7][25] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\ann.ReLU_out[8][9] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\ann.ReLU_out[3][23] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\ann.ReLU_out[7][24] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\ann.ReLU_out[9][8] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\ann.ReLU_out[5][8] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\ann.ReLU_out[2][26] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\ann.ReLU_out[1][23] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\ann.ReLU_out[1][26] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0152_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\ann.ReLU_out[9][9] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\ann.ReLU_out[8][11] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\ann.ReLU_out[1][24] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\ann.ReLU_out[2][24] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\ann.ReLU_out[4][24] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\ann.ReLU_out[4][17] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\ann.ReLU_out[5][16] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\ann.ReLU_out[1][19] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\ann.ReLU_out[8][10] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\ann.ReLU_out[7][12] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\ann.ReLU_out[0][29] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\ann.ReLU_out[4][6] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\ann.ReLU_out[3][1] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\ann.ReLU_out[6][24] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\ann.ReLU_out[5][24] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\ann.ReLU_out[3][29] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\ann.ReLU_out[9][1] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\ann.ReLU_out[2][6] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\ann.ReLU_out[4][21] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\ann.ReLU_out[9][16] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\ann.ReLU_out[9][23] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0156_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0164_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\ann.ReLU_out[3][25] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\ann.ReLU_out[8][26] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\ann.ReLU_out[1][17] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\ann.in_ff[2][1] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\ann.ReLU_out[7][11] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\ann.ReLU_out[6][1] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\ann.ReLU_out[7][6] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\ann.ReLU_out[1][25] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\ann.ReLU_out[9][28] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\ann.ReLU_out[6][18] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\ann.ReLU_out[0][10] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\ann.ReLU_out[8][16] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\ann.ReLU_out[3][22] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\ann.ReLU_out[5][6] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0296_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\ann.ReLU_out[4][22] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\ann.ReLU_out[7][9] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\ann.ReLU_out[2][23] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\ann.ReLU_out[2][22] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\ann.ReLU_out[3][12] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\ann.ReLU_out[9][11] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0145_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\ann.ReLU_out[4][26] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\ann.ReLU_out[6][21] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\ann.ReLU_out[3][6] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\ann.ReLU_out[9][6] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\ann.ReLU_out[8][22] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\ann.ReLU_out[2][9] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\ann.ReLU_out[5][23] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\ann.ReLU_out[6][27] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\ann.ReLU_out[9][3] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\ann.ReLU_out[7][22] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\ann.ReLU_out[0][7] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\ann.ReLU_out[6][11] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\ann.ReLU_out[4][23] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\ann.ReLU_out[6][6] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\ann.ReLU_out[6][26] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\ann.ReLU_out[6][9] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\ann.ReLU_out[2][8] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\ann.ReLU_out[8][12] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\ann.ReLU_out[3][18] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\ann.ReLU_out[8][4] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\ann.ReLU_out[6][23] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0142_),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\ann.ReLU_out[4][1] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\ann.ReLU_out[3][17] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\ann.ReLU_out[1][14] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\ann.ReLU_out[7][8] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\ann.ReLU_out[6][29] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\ann.ReLU_out[2][13] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\ann.ReLU_out[3][2] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\ann.ReLU_out[7][26] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\ann.ReLU_out[3][3] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\ann.ReLU_out[2][1] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\ann.ReLU_out[0][16] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\ann.ReLU_out[2][12] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\ann.ReLU_out[4][29] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\ann.ReLU_out[5][12] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\ann.ReLU_out[2][30] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\ann.ReLU_out[7][10] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\ann.ReLU_out[7][5] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\ann.ReLU_out[9][10] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\ann.ReLU_out[7][1] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\ann.ReLU_out[3][4] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\ann.ReLU_out[8][2] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0151_),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\ann.ReLU_out[7][2] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\ann.ReLU_out[3][16] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\ann.ReLU_out[7][4] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\ann.ReLU_out[8][25] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\ann.ReLU_out[5][2] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\ann.ReLU_out[8][13] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\ann.ReLU_out[1][2] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\ann.ReLU_out[2][14] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\ann.ReLU_out[1][6] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\ann.ReLU_out[3][7] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\ann.ReLU_out[0][23] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\ann.ReLU_out[5][4] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\ann.ReLU_out[2][2] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\ann.ReLU_out[5][1] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\ann.ReLU_out[5][17] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\ann.ReLU_out[3][14] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\ann.ReLU_out[6][25] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\ann.ReLU_out[6][5] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\ann.ReLU_out[2][4] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\ann.ReLU_out[2][5] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\ann.ReLU_out[8][7] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0158_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\ann.ReLU_out[5][26] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\ann.ReLU_out[3][5] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\ann.ReLU_out[4][2] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\ann.ReLU_out[1][5] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\ann.ReLU_out[7][16] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\ann.ReLU_out[5][20] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\ann.ReLU_out[1][3] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\ann.ReLU_out[4][4] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\ann.ReLU_out[6][4] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\ann.ReLU_out[6][2] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\ann.ReLU_out[0][2] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\ann.ReLU_out[2][3] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\ann.ReLU_out[8][8] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\ann.ReLU_out[3][13] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\ann.ReLU_out[2][11] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\ann.ReLU_out[9][24] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\ann.ReLU_out[9][5] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\ann.ReLU_out[8][5] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\ann.ReLU_out[2][7] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\ann.ReLU_out[4][5] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\ann.ReLU_out[5][9] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\ann.ReLU_out[0][30] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0137_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\ann.ReLU_out[7][3] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\ann.ReLU_out[5][7] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\ann.ReLU_out[1][9] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\ann.ReLU_out[5][21] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\ann.ReLU_out[4][12] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\ann.ReLU_out[5][30] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\ann.ReLU_out[8][3] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\ann.ReLU_out[1][7] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\ann.ReLU_out[5][5] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\ann.ReLU_out[5][10] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\ann.ReLU_out[0][20] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\ann.ReLU_out[7][7] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\ann.ReLU_out[4][3] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\ann.ReLU_out[1][4] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\ann.ReLU_out[3][11] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\ann.ReLU_out[6][28] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\ann.ReLU_out[5][11] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\ann.ReLU_out[5][3] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\ann.ReLU_out[4][13] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\ann.ReLU_out[4][7] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\ann.ReLU_out[1][1] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0155_),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\ann.ReLU_out[6][3] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\ann.ReLU_out[7][13] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\ann.ReLU_out[9][7] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\ann.ReLU_out[9][2] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\ann.ReLU_out[6][7] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\ann.ReLU_out[2][10] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\ann.ReLU_out[8][6] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\ann.ReLU_out[9][26] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\ann.ReLU_out[3][9] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\ann.ReLU_out[8][14] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\ann.ReLU_out[0][0] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\ann.in_ff[2][0] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\ann.ReLU_out[4][11] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\ann.ReLU_out[8][28] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\ann.ReLU_out[8][17] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\ann.ReLU_out[6][14] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\ann.ReLU_out[4][20] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\ann.ReLU_out[3][20] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\ann.ReLU_out[4][9] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\ann.ReLU_out[7][14] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\ann.ReLU_out[7][28] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0135_),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\ann.ReLU_out[1][11] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\ann.ReLU_out[5][13] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\ann.ReLU_out[4][10] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\ann.ReLU_out[1][28] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\ann.ReLU_out[2][18] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\ann.ReLU_out[9][21] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\ann.ReLU_out[3][21] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\ann.ReLU_out[5][14] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\ann.ReLU_out[1][13] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\ann.ReLU_out[4][18] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\ann.ReLU_out[0][24] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\ann.ReLU_out[1][12] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\ann.ReLU_out[3][10] ),
    .X(net605));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold352 (.A(\ann.ReLU_out[9][4] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\ann.ReLU_out[1][20] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\ann.ReLU_out[9][25] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\ann.ReLU_out[5][28] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\ann.ReLU_out[8][30] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\ann.in_ff[2][12] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\ann.ReLU_out[2][27] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\ann.ReLU_out[7][30] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0159_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\ann.ReLU_out[6][13] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\ann.ReLU_out[5][18] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\ann.ReLU_out[4][14] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\ann.ReLU_out[9][14] ),
    .X(net617));
 sky130_fd_sc_hd__buf_1 hold364 (.A(net790),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\ann.in_ff[2][7] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\ann.ReLU_out[9][12] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\ann.ReLU_out[2][20] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\ann.ReLU_out[4][25] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\ann.ReLU_out[4][30] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\ann.ReLU_out[0][6] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\ann.ReLU_out[5][27] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\ann.in_ff[2][4] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\ann.ReLU_out[3][26] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\ann.ReLU_out[7][27] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\ann.ReLU_out[4][27] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\ann.ReLU_out[5][19] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\ann.in_ff[2][6] ),
    .X(net630));
 sky130_fd_sc_hd__buf_1 hold377 (.A(\ann.ReLU_out[9][30] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\ann.ReLU_out[8][21] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\ann.ReLU_out[7][21] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0141_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\ann.ReLU_out[8][20] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\ann.in_ff[2][5] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\ann.ReLU_out[9][18] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\ann.ReLU_out[7][17] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\ann.ReLU_out[1][10] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\ann.ReLU_out[2][21] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\ann.ReLU_out[7][29] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\ann.ReLU_out[7][19] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\ann.in_ff[2][8] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\ann.ReLU_out[8][27] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\ann.ReLU_out[0][27] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\ann.temp[24] ),
    .X(net644));
 sky130_fd_sc_hd__buf_1 hold391 (.A(net791),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\ann.ReLU_out[8][19] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\ann.ReLU_out[1][29] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\ann.ReLU_out[1][21] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\ann.in_ff[2][11] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\ann.ReLU_out[9][13] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\ann.ReLU_out[6][20] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\ann.in_ff[2][2] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\ann.in_ff[2][3] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0165_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0162_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\ann.in_ff[2][15] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\ann.ReLU_out[6][19] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\ann.temp[25] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\ann.ReLU_out[9][22] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\ann.temp[23] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\ann.ReLU_out[9][20] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\ann.in_ff[2][9] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\ann.in_ff[2][13] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\ann.in_ff[2][14] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\ann.ReLU_out[7][20] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\ann.ReLU_out[0][4] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\ann.ReLU_out[9][27] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\ann.ReLU_out[1][27] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\ann.temp[20] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\ann.ReLU_out[3][15] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\ann.in_ff[2][10] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\ann.ReLU_out[8][15] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\ann.ReLU_out[2][19] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\ann.ReLU_out[1][15] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\ann.ReLU_out[9][29] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\ann.ReLU_out[9][19] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0139_),
    .X(net296));
 sky130_fd_sc_hd__buf_1 hold420 (.A(net792),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\ann.temp[21] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\ann.ReLU_out[8][29] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\ann.ReLU_out[6][15] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\ann.ReLU_out[2][25] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\ann.ReLU_out[7][18] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\ann.in_ff[0][0] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\ann.ReLU_out[5][15] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\ann.ReLU_out[9][15] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\ann.in_ff[0][1] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\ann.ReLU_out[0][5] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\ann.ReLU_out[4][15] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\ann.in_ff[0][9] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\ann.in_ff[0][3] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\ann.ReLU_out[7][15] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\ann.in_ff[0][2] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\ann.in_ff[0][7] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\ann.in_ff[0][6] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\ann.ReLU_out[4][19] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\ann.in_ff[0][4] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\ann.in_ff[0][8] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0140_),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\ann.in_ff[0][5] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\ann.ReLU_out[2][15] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\ann.in_ff[0][14] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\ann.ReLU_out[1][30] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\ann.in_ff[0][11] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\ann.in_ff[0][10] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\ann.in_ff[0][12] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\ann.ReLU_out[5][25] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\ann.X[31] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\ann.in_ff[0][15] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\ann.ReLU_out[0][22] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\ann.bias[18] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\ann.X[28] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\ann.in_ff[0][13] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\ann.ReLU_out[3][27] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\ann.ReLU_out[8][18] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\ann.bias[9] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\ann.bias[6] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\ann.bias[21] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\ann.temp[15] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\ann.X[29] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0157_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\ann.X[18] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\ann.X[10] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\ann.X[30] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\ann.temp[29] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\ann.X[0] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\ann.X[15] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\ann.X[4] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\ann.X[17] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\ann.X[26] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\ann.X[9] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\ann.ReLU_out[0][11] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\ann.bias[19] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\ann.bias[3] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\ann.X[23] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\ann.bias[12] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\ann.ReLU_out[3][19] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\ann.X[3] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\ann.bias[7] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\ann.state[0] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\ann.bias[11] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\ann.X[8] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0146_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\ann.bias[20] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\ann.bias[31] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\ann.X[1] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\ann.X[2] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\ann.X[19] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\ann.X[7] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\ann.bias[28] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\ann.X[16] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\ann.bias[30] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\ann.temp[28] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\ann.ReLU_out[0][3] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\ann.bias[10] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\ann.bias[1] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\ann.X[14] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\ann.temp[9] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\ann.ReLU_out[1][22] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\ann.bias[15] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\ann.temp[10] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\ann.X[22] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\ann.X[12] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\ann.temp[11] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\ann.ReLU_out[0][14] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0138_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\ann.bias[17] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\ann.temp[16] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\ann.X[27] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\ann.temp[27] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\ann.temp[8] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\ann.bias[2] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\ann.bias[8] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\ann.bias[4] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\ann.bias[23] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\ann.X[6] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\ann.ReLU_out[0][8] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\ann.bias[5] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\ann.temp[17] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\ann.X[13] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\ann.X[11] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\ann.X[20] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\ann.X[24] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\ann.bias[22] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\ann.bias[13] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\ann.bias[14] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\ann.temp[26] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0143_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\ann.temp[19] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\ann.bias[25] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\ann.X[25] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\ann.X[21] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\ann.bias[0] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\ann.bias[24] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\ann.bias[29] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\ann.X[5] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\ann.temp[18] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\ann.bias[16] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\ann.ReLU_out[0][19] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\ann.temp[30] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\ann.temp[22] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\ann.bias[26] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\ann.bias[27] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\ann.temp[30] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\ann.state[0] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\ann.ReLU_out[2][28] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\ann.ReLU_out[3][28] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\ann.ReLU_out[4][28] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0154_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\ann.ReLU_out[0][25] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0160_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\ann.ReLU_out[0][28] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0163_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\ann.temp[14] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0149_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0118_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\ann.temp[13] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0117_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\ann.ReLU_out[0][15] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0150_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\ann.ReLU_out[0][26] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0161_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\ann.ReLU_out[6][30] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0351_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\ann.ReLU_out[1][0] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\ann.ReLU_out[0][9] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0166_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\ann.ReLU_out[2][0] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0197_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\ann.in_ff[1][7] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0532_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\ann.temp[5] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0109_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\ann.in_ff[1][0] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0525_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\ann.temp[7] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0144_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0111_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\ann.ReLU_out[6][17] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0338_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\ann.ReLU_out[6][8] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0329_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\ann.temp[12] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0116_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\ann.ReLU_out[3][0] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0228_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\ann.temp[2] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\ann.ReLU_out[0][1] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0106_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\ann.in_ff[1][1] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0526_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\ann.ReLU_out[5][0] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0290_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\ann.temp[3] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0107_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\ann.temp[4] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0108_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\ann.temp[0] ),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(io_in[10]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_16 input10 (.A(io_in[19]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 input11 (.A(io_in[20]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 input12 (.A(io_in[21]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input13 (.A(io_in[22]),
    .X(net13));
 sky130_fd_sc_hd__buf_8 input14 (.A(io_in[23]),
    .X(net14));
 sky130_fd_sc_hd__buf_8 input15 (.A(io_in[24]),
    .X(net15));
 sky130_fd_sc_hd__buf_8 input16 (.A(io_in[25]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_8 input17 (.A(io_in[26]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_8 input18 (.A(io_in[27]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(io_in[28]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(io_in[11]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(io_in[29]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(io_in[30]),
    .X(net21));
 sky130_fd_sc_hd__buf_8 input22 (.A(io_in[31]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 input23 (.A(io_in[32]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(io_in[33]),
    .X(net24));
 sky130_fd_sc_hd__buf_8 input25 (.A(io_in[35]),
    .X(net25));
 sky130_fd_sc_hd__buf_8 input26 (.A(io_in[36]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_16 input27 (.A(io_in[37]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(io_in[7]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_8 input29 (.A(io_in[8]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(io_in[12]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input30 (.A(io_in[9]),
    .X(net30));
 sky130_fd_sc_hd__buf_12 input31 (.A(wb_rst_i),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(io_in[13]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(io_in[14]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(io_in[15]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(io_in[16]),
    .X(net7));
 sky130_fd_sc_hd__buf_8 input8 (.A(io_in[17]),
    .X(net8));
 sky130_fd_sc_hd__buf_8 input9 (.A(io_in[18]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 max_cap57 (.A(_1972_),
    .X(net57));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(io_out[6]));
 sky130_fd_sc_hd__conb_1 user_proj_example_219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 user_proj_example_220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 user_proj_example_221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 user_proj_example_222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 user_proj_example_224 (.HI(net224));
 sky130_fd_sc_hd__conb_1 user_proj_example_225 (.HI(net225));
 sky130_fd_sc_hd__conb_1 user_proj_example_226 (.HI(net226));
 sky130_fd_sc_hd__conb_1 user_proj_example_227 (.HI(net227));
 sky130_fd_sc_hd__conb_1 user_proj_example_228 (.HI(net228));
 sky130_fd_sc_hd__conb_1 user_proj_example_229 (.HI(net229));
 sky130_fd_sc_hd__conb_1 user_proj_example_230 (.HI(net230));
 sky130_fd_sc_hd__conb_1 user_proj_example_231 (.HI(net231));
 sky130_fd_sc_hd__conb_1 user_proj_example_232 (.HI(net232));
 sky130_fd_sc_hd__conb_1 user_proj_example_233 (.HI(net233));
 sky130_fd_sc_hd__conb_1 user_proj_example_234 (.HI(net234));
 sky130_fd_sc_hd__conb_1 user_proj_example_235 (.HI(net235));
 sky130_fd_sc_hd__conb_1 user_proj_example_236 (.HI(net236));
 sky130_fd_sc_hd__conb_1 user_proj_example_237 (.HI(net237));
 sky130_fd_sc_hd__conb_1 user_proj_example_238 (.HI(net238));
 sky130_fd_sc_hd__conb_1 user_proj_example_239 (.HI(net239));
 sky130_fd_sc_hd__conb_1 user_proj_example_240 (.HI(net240));
 sky130_fd_sc_hd__conb_1 user_proj_example_241 (.HI(net241));
 sky130_fd_sc_hd__conb_1 user_proj_example_242 (.HI(net242));
 sky130_fd_sc_hd__conb_1 user_proj_example_243 (.HI(net243));
 sky130_fd_sc_hd__conb_1 user_proj_example_244 (.HI(net244));
 sky130_fd_sc_hd__conb_1 user_proj_example_245 (.HI(net245));
 sky130_fd_sc_hd__conb_1 user_proj_example_246 (.HI(net246));
 sky130_fd_sc_hd__conb_1 user_proj_example_247 (.HI(net247));
 sky130_fd_sc_hd__conb_1 user_proj_example_248 (.HI(net248));
 sky130_fd_sc_hd__conb_1 user_proj_example_249 (.HI(net249));
 sky130_fd_sc_hd__conb_1 user_proj_example_250 (.HI(net250));
 sky130_fd_sc_hd__conb_1 user_proj_example_251 (.HI(net251));
 sky130_fd_sc_hd__conb_1 user_proj_example_252 (.HI(net252));
 sky130_fd_sc_hd__conb_1 user_proj_example_253 (.HI(net253));
 sky130_fd_sc_hd__conb_1 user_proj_example_254 (.HI(net254));
 assign io_oeb[10] = net227;
 assign io_oeb[11] = net228;
 assign io_oeb[12] = net229;
 assign io_oeb[13] = net230;
 assign io_oeb[14] = net231;
 assign io_oeb[15] = net232;
 assign io_oeb[16] = net233;
 assign io_oeb[17] = net234;
 assign io_oeb[18] = net235;
 assign io_oeb[19] = net236;
 assign io_oeb[20] = net237;
 assign io_oeb[21] = net238;
 assign io_oeb[22] = net239;
 assign io_oeb[23] = net240;
 assign io_oeb[24] = net241;
 assign io_oeb[25] = net242;
 assign io_oeb[26] = net243;
 assign io_oeb[27] = net244;
 assign io_oeb[28] = net245;
 assign io_oeb[29] = net246;
 assign io_oeb[30] = net247;
 assign io_oeb[31] = net248;
 assign io_oeb[32] = net249;
 assign io_oeb[33] = net250;
 assign io_oeb[34] = net251;
 assign io_oeb[35] = net252;
 assign io_oeb[36] = net253;
 assign io_oeb[37] = net254;
 assign io_oeb[3] = net219;
 assign io_oeb[4] = net220;
 assign io_oeb[5] = net221;
 assign io_oeb[6] = net222;
 assign io_oeb[7] = net224;
 assign io_oeb[8] = net225;
 assign io_oeb[9] = net226;
endmodule

