magic
tech sky130A
magscale 1 2
timestamp 1702347434
<< obsli1 >>
rect 1104 2159 38824 597329
<< obsm1 >>
rect 934 2128 39086 597360
<< metal2 >>
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 938 856 39080 597349
rect 938 800 9898 856
rect 10066 800 29862 856
rect 30030 800 39080 856
<< metal3 >>
rect 39200 590248 40000 590368
rect 0 586984 800 587104
rect 39200 573656 40000 573776
rect 0 569576 800 569696
rect 39200 557064 40000 557184
rect 0 552168 800 552288
rect 39200 540472 40000 540592
rect 0 534760 800 534880
rect 39200 523880 40000 524000
rect 0 517352 800 517472
rect 39200 507288 40000 507408
rect 0 499944 800 500064
rect 39200 490696 40000 490816
rect 0 482536 800 482656
rect 39200 474104 40000 474224
rect 0 465128 800 465248
rect 39200 457512 40000 457632
rect 0 447720 800 447840
rect 39200 440920 40000 441040
rect 0 430312 800 430432
rect 39200 424328 40000 424448
rect 0 412904 800 413024
rect 39200 407736 40000 407856
rect 0 395496 800 395616
rect 39200 391144 40000 391264
rect 0 378088 800 378208
rect 39200 374552 40000 374672
rect 0 360680 800 360800
rect 39200 357960 40000 358080
rect 0 343272 800 343392
rect 39200 341368 40000 341488
rect 0 325864 800 325984
rect 39200 324776 40000 324896
rect 0 308456 800 308576
rect 39200 308184 40000 308304
rect 39200 291592 40000 291712
rect 0 291048 800 291168
rect 39200 275000 40000 275120
rect 0 273640 800 273760
rect 39200 258408 40000 258528
rect 0 256232 800 256352
rect 39200 241816 40000 241936
rect 0 238824 800 238944
rect 39200 225224 40000 225344
rect 0 221416 800 221536
rect 39200 208632 40000 208752
rect 0 204008 800 204128
rect 39200 192040 40000 192160
rect 0 186600 800 186720
rect 39200 175448 40000 175568
rect 0 169192 800 169312
rect 39200 158856 40000 158976
rect 0 151784 800 151904
rect 39200 142264 40000 142384
rect 0 134376 800 134496
rect 39200 125672 40000 125792
rect 0 116968 800 117088
rect 39200 109080 40000 109200
rect 0 99560 800 99680
rect 39200 92488 40000 92608
rect 0 82152 800 82272
rect 39200 75896 40000 76016
rect 0 64744 800 64864
rect 39200 59304 40000 59424
rect 0 47336 800 47456
rect 39200 42712 40000 42832
rect 0 29928 800 30048
rect 39200 26120 40000 26240
rect 0 12520 800 12640
rect 39200 9528 40000 9648
<< obsm3 >>
rect 798 590448 39200 597345
rect 798 590168 39120 590448
rect 798 587184 39200 590168
rect 880 586904 39200 587184
rect 798 573856 39200 586904
rect 798 573576 39120 573856
rect 798 569776 39200 573576
rect 880 569496 39200 569776
rect 798 557264 39200 569496
rect 798 556984 39120 557264
rect 798 552368 39200 556984
rect 880 552088 39200 552368
rect 798 540672 39200 552088
rect 798 540392 39120 540672
rect 798 534960 39200 540392
rect 880 534680 39200 534960
rect 798 524080 39200 534680
rect 798 523800 39120 524080
rect 798 517552 39200 523800
rect 880 517272 39200 517552
rect 798 507488 39200 517272
rect 798 507208 39120 507488
rect 798 500144 39200 507208
rect 880 499864 39200 500144
rect 798 490896 39200 499864
rect 798 490616 39120 490896
rect 798 482736 39200 490616
rect 880 482456 39200 482736
rect 798 474304 39200 482456
rect 798 474024 39120 474304
rect 798 465328 39200 474024
rect 880 465048 39200 465328
rect 798 457712 39200 465048
rect 798 457432 39120 457712
rect 798 447920 39200 457432
rect 880 447640 39200 447920
rect 798 441120 39200 447640
rect 798 440840 39120 441120
rect 798 430512 39200 440840
rect 880 430232 39200 430512
rect 798 424528 39200 430232
rect 798 424248 39120 424528
rect 798 413104 39200 424248
rect 880 412824 39200 413104
rect 798 407936 39200 412824
rect 798 407656 39120 407936
rect 798 395696 39200 407656
rect 880 395416 39200 395696
rect 798 391344 39200 395416
rect 798 391064 39120 391344
rect 798 378288 39200 391064
rect 880 378008 39200 378288
rect 798 374752 39200 378008
rect 798 374472 39120 374752
rect 798 360880 39200 374472
rect 880 360600 39200 360880
rect 798 358160 39200 360600
rect 798 357880 39120 358160
rect 798 343472 39200 357880
rect 880 343192 39200 343472
rect 798 341568 39200 343192
rect 798 341288 39120 341568
rect 798 326064 39200 341288
rect 880 325784 39200 326064
rect 798 324976 39200 325784
rect 798 324696 39120 324976
rect 798 308656 39200 324696
rect 880 308384 39200 308656
rect 880 308376 39120 308384
rect 798 308104 39120 308376
rect 798 291792 39200 308104
rect 798 291512 39120 291792
rect 798 291248 39200 291512
rect 880 290968 39200 291248
rect 798 275200 39200 290968
rect 798 274920 39120 275200
rect 798 273840 39200 274920
rect 880 273560 39200 273840
rect 798 258608 39200 273560
rect 798 258328 39120 258608
rect 798 256432 39200 258328
rect 880 256152 39200 256432
rect 798 242016 39200 256152
rect 798 241736 39120 242016
rect 798 239024 39200 241736
rect 880 238744 39200 239024
rect 798 225424 39200 238744
rect 798 225144 39120 225424
rect 798 221616 39200 225144
rect 880 221336 39200 221616
rect 798 208832 39200 221336
rect 798 208552 39120 208832
rect 798 204208 39200 208552
rect 880 203928 39200 204208
rect 798 192240 39200 203928
rect 798 191960 39120 192240
rect 798 186800 39200 191960
rect 880 186520 39200 186800
rect 798 175648 39200 186520
rect 798 175368 39120 175648
rect 798 169392 39200 175368
rect 880 169112 39200 169392
rect 798 159056 39200 169112
rect 798 158776 39120 159056
rect 798 151984 39200 158776
rect 880 151704 39200 151984
rect 798 142464 39200 151704
rect 798 142184 39120 142464
rect 798 134576 39200 142184
rect 880 134296 39200 134576
rect 798 125872 39200 134296
rect 798 125592 39120 125872
rect 798 117168 39200 125592
rect 880 116888 39200 117168
rect 798 109280 39200 116888
rect 798 109000 39120 109280
rect 798 99760 39200 109000
rect 880 99480 39200 99760
rect 798 92688 39200 99480
rect 798 92408 39120 92688
rect 798 82352 39200 92408
rect 880 82072 39200 82352
rect 798 76096 39200 82072
rect 798 75816 39120 76096
rect 798 64944 39200 75816
rect 880 64664 39200 64944
rect 798 59504 39200 64664
rect 798 59224 39120 59504
rect 798 47536 39200 59224
rect 880 47256 39200 47536
rect 798 42912 39200 47256
rect 798 42632 39120 42912
rect 798 30128 39200 42632
rect 880 29848 39200 30128
rect 798 26320 39200 29848
rect 798 26040 39120 26320
rect 798 12720 39200 26040
rect 880 12440 39200 12720
rect 798 9728 39200 12440
rect 798 9448 39120 9728
rect 798 2143 39200 9448
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
<< obsm4 >>
rect 1715 77147 4128 438157
rect 4608 77147 19488 438157
rect 19968 77147 34848 438157
rect 35328 77147 36741 438157
<< labels >>
rlabel metal3 s 39200 241816 40000 241936 6 io_in[10]
port 1 nsew signal input
rlabel metal3 s 39200 275000 40000 275120 6 io_in[11]
port 2 nsew signal input
rlabel metal3 s 39200 308184 40000 308304 6 io_in[12]
port 3 nsew signal input
rlabel metal3 s 39200 341368 40000 341488 6 io_in[13]
port 4 nsew signal input
rlabel metal3 s 39200 374552 40000 374672 6 io_in[14]
port 5 nsew signal input
rlabel metal3 s 39200 407736 40000 407856 6 io_in[15]
port 6 nsew signal input
rlabel metal3 s 39200 440920 40000 441040 6 io_in[16]
port 7 nsew signal input
rlabel metal3 s 39200 474104 40000 474224 6 io_in[17]
port 8 nsew signal input
rlabel metal3 s 39200 507288 40000 507408 6 io_in[18]
port 9 nsew signal input
rlabel metal3 s 39200 540472 40000 540592 6 io_in[19]
port 10 nsew signal input
rlabel metal3 s 39200 573656 40000 573776 6 io_in[20]
port 11 nsew signal input
rlabel metal3 s 0 586984 800 587104 6 io_in[21]
port 12 nsew signal input
rlabel metal3 s 0 552168 800 552288 6 io_in[22]
port 13 nsew signal input
rlabel metal3 s 0 517352 800 517472 6 io_in[23]
port 14 nsew signal input
rlabel metal3 s 0 482536 800 482656 6 io_in[24]
port 15 nsew signal input
rlabel metal3 s 0 447720 800 447840 6 io_in[25]
port 16 nsew signal input
rlabel metal3 s 0 412904 800 413024 6 io_in[26]
port 17 nsew signal input
rlabel metal3 s 0 378088 800 378208 6 io_in[27]
port 18 nsew signal input
rlabel metal3 s 0 343272 800 343392 6 io_in[28]
port 19 nsew signal input
rlabel metal3 s 0 308456 800 308576 6 io_in[29]
port 20 nsew signal input
rlabel metal3 s 0 273640 800 273760 6 io_in[30]
port 21 nsew signal input
rlabel metal3 s 0 238824 800 238944 6 io_in[31]
port 22 nsew signal input
rlabel metal3 s 0 204008 800 204128 6 io_in[32]
port 23 nsew signal input
rlabel metal3 s 0 169192 800 169312 6 io_in[33]
port 24 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 io_in[34]
port 25 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 io_in[35]
port 26 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_in[36]
port 27 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 io_in[37]
port 28 nsew signal input
rlabel metal3 s 39200 142264 40000 142384 6 io_in[7]
port 29 nsew signal input
rlabel metal3 s 39200 175448 40000 175568 6 io_in[8]
port 30 nsew signal input
rlabel metal3 s 39200 208632 40000 208752 6 io_in[9]
port 31 nsew signal input
rlabel metal3 s 39200 258408 40000 258528 6 io_oeb[10]
port 32 nsew signal output
rlabel metal3 s 39200 291592 40000 291712 6 io_oeb[11]
port 33 nsew signal output
rlabel metal3 s 39200 324776 40000 324896 6 io_oeb[12]
port 34 nsew signal output
rlabel metal3 s 39200 357960 40000 358080 6 io_oeb[13]
port 35 nsew signal output
rlabel metal3 s 39200 391144 40000 391264 6 io_oeb[14]
port 36 nsew signal output
rlabel metal3 s 39200 424328 40000 424448 6 io_oeb[15]
port 37 nsew signal output
rlabel metal3 s 39200 457512 40000 457632 6 io_oeb[16]
port 38 nsew signal output
rlabel metal3 s 39200 490696 40000 490816 6 io_oeb[17]
port 39 nsew signal output
rlabel metal3 s 39200 523880 40000 524000 6 io_oeb[18]
port 40 nsew signal output
rlabel metal3 s 39200 557064 40000 557184 6 io_oeb[19]
port 41 nsew signal output
rlabel metal3 s 39200 590248 40000 590368 6 io_oeb[20]
port 42 nsew signal output
rlabel metal3 s 0 569576 800 569696 6 io_oeb[21]
port 43 nsew signal output
rlabel metal3 s 0 534760 800 534880 6 io_oeb[22]
port 44 nsew signal output
rlabel metal3 s 0 499944 800 500064 6 io_oeb[23]
port 45 nsew signal output
rlabel metal3 s 0 465128 800 465248 6 io_oeb[24]
port 46 nsew signal output
rlabel metal3 s 0 430312 800 430432 6 io_oeb[25]
port 47 nsew signal output
rlabel metal3 s 0 395496 800 395616 6 io_oeb[26]
port 48 nsew signal output
rlabel metal3 s 0 360680 800 360800 6 io_oeb[27]
port 49 nsew signal output
rlabel metal3 s 0 325864 800 325984 6 io_oeb[28]
port 50 nsew signal output
rlabel metal3 s 0 291048 800 291168 6 io_oeb[29]
port 51 nsew signal output
rlabel metal3 s 0 256232 800 256352 6 io_oeb[30]
port 52 nsew signal output
rlabel metal3 s 0 221416 800 221536 6 io_oeb[31]
port 53 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 io_oeb[32]
port 54 nsew signal output
rlabel metal3 s 0 151784 800 151904 6 io_oeb[33]
port 55 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 io_oeb[34]
port 56 nsew signal output
rlabel metal3 s 0 82152 800 82272 6 io_oeb[35]
port 57 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 io_oeb[36]
port 58 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 io_oeb[37]
port 59 nsew signal output
rlabel metal3 s 39200 26120 40000 26240 6 io_oeb[3]
port 60 nsew signal output
rlabel metal3 s 39200 59304 40000 59424 6 io_oeb[4]
port 61 nsew signal output
rlabel metal3 s 39200 92488 40000 92608 6 io_oeb[5]
port 62 nsew signal output
rlabel metal3 s 39200 125672 40000 125792 6 io_oeb[6]
port 63 nsew signal output
rlabel metal3 s 39200 158856 40000 158976 6 io_oeb[7]
port 64 nsew signal output
rlabel metal3 s 39200 192040 40000 192160 6 io_oeb[8]
port 65 nsew signal output
rlabel metal3 s 39200 225224 40000 225344 6 io_oeb[9]
port 66 nsew signal output
rlabel metal3 s 39200 9528 40000 9648 6 io_out[3]
port 67 nsew signal output
rlabel metal3 s 39200 42712 40000 42832 6 io_out[4]
port 68 nsew signal output
rlabel metal3 s 39200 75896 40000 76016 6 io_out[5]
port 69 nsew signal output
rlabel metal3 s 39200 109080 40000 109200 6 io_out[6]
port 70 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 71 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 71 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 72 nsew ground bidirectional
rlabel metal2 s 9954 0 10010 800 6 wb_clk_i
port 73 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_rst_i
port 74 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 21615572
string GDS_FILE /home/paras22167/Caravel/caravel_user_project/openlane/user_proj_example/runs/23_12_12_07_36/results/signoff/user_proj_example.magic.gds
string GDS_START 1035094
<< end >>

